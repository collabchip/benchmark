module pci_bridge32 (
x13786,
x13626,
x12891,
x6501,
x4455,
x13353,
x13185,
x4489,
x13674,
x13779,
x13712,
x5001,
x13364,
x4851,
x4420,
x4295,
x13520,
x4886,
x13156,
x13808,
x4932,
x13134,
x13058,
x4743,
x13069,
x4701,
x12902,
x13698,
x13567,
x13038,
x4392,
x4861,
x4496,
x4821,
x192485,
x13004,
x12780,
x13994,
x4778,
x4635,
x13330,
x4323,
x12969,
x13560,
x13031,
x13750,
x12922,
x13252,
x4576,
x13018,
x13047,
x13494,
x13208,
x13174,
x13433,
x13594,
x13440,
x13126,
x13403,
x4805,
x13193,
x13474,
x13341,
x13423,
x13612,
x13843,
x13100,
x13663,
x12843,
x13234,
x13633,
x4764,
x12810,
x12991,
x13011,
x13541,
x13025,
x13396,
x4707,
x13291,
x13644,
x13447,
x13654,
x13093,
x4964,
x13414,
x4840,
x13145,
x13263,
x12929,
x13733,
x13853,
x4812,
x13547,
x13576,
x13921,
x12915,
x13553,
x4771,
x12962,
x13514,
x4733,
x13605,
x13271,
x13863,
x4347,
x4919,
x13742,
x192486,
x13534,
x13833,
x13501,
x14005,
x13722,
x13761,
x13508,
x13684,
x13705,
x4538,
x13527,
x13969,
x13884,
x13797,
x4796,
x13586,
x4367,
x13950,
x4831,
x13984,
x12940,
x4570,
x12980,
x13385,
x13482,
x13619,
x13464,
x4869,
x4514,
x13115,
x13772,
x4448,
x13488,
x12768,
x4503,
x4902,
x12955,
x4788,
x4693,
x13374,
x192484,
x4607,
x13086,
x13826,
x13815,
x4757,
x13077,
x13457,
x4561,
x13163,
x13870,
x4254,
x4667,
x757,
x749,
x291,
x508,
x971,
x2633,
x729,
x4227,
x4234,
x451,
x1244,
x815,
x3122,
x1087,
x3996,
x1032,
x912,
x4059,
x1024,
x3954,
x3524,
x2693,
x468,
x378,
x1215,
x225,
x364,
x3816,
x852,
x594,
x1721,
x712,
x2981,
x1745,
x879,
x1062,
x352,
x3372,
x420,
x1575,
x4214,
x4023,
x827,
x753,
x764,
x697,
x521,
x3028,
x9,
x4192,
x3803,
x3762,
x170,
x186,
x3861,
x240,
x845,
x725,
x4154,
x926,
x4049,
x132,
x2594,
x1152,
x871,
x3258,
x338,
x3968,
x2805,
x863,
x434,
x1885,
x3561,
x963,
x4082,
x52,
x20,
x4115,
x2068,
x1039,
x1778,
x3925,
x2542,
x1340,
x808,
x0,
x2308,
x1977,
x3418,
x3604,
x27,
x1855,
x2494,
x2006,
x4143,
x2100,
x4104,
x2856,
x890,
x1804,
x2451,
x3904,
x3847,
x3712,
x608,
x1829,
x1174,
x1532,
x1383,
x3485,
x76,
x771,
x831,
x4070,
x683,
x820,
x1639,
x1690,
x2746,
x306,
x2908,
x2400,
x778,
x3938,
x999,
x3830,
x3685,
x3874,
x480,
x956,
x105,
x1597,
x2169,
x801,
x3451,
x2355,
x933,
x735,
x4093,
x649,
x1912,
x641,
x919,
x661,
x653,
x2230,
x3156,
x1070,
x1130,
x2261,
x552,
x677,
x494,
x905,
x3327,
x1195,
x785,
x1305,
x2948,
x43,
x719,
x668,
x838,
x4132,
x4011,
x742,
x154,
x1016,
x690,
x703,
x4036,
x563,
x2041,
x886,
x1010,
x34,
x394,
x1281,
x4166,
x3207,
x2133,
x3079,
x898,
x1500,
x258,
x324,
x3288,
x789,
x275,
x1935,
x1467,
x3891,
x208,
x406,
x577,
x1107,
x1667,
x1428,
x794,
x626,
x2195,
x4204,
x856,
x4179,
x3651,
x3983,
x534);

// Start PIs
input x13786;
input x13626;
input x12891;
input x6501;
input x4455;
input x13353;
input x13185;
input x4489;
input x13674;
input x13779;
input x13712;
input x5001;
input x13364;
input x4851;
input x4420;
input x4295;
input x13520;
input x4886;
input x13156;
input x13808;
input x4932;
input x13134;
input x13058;
input x4743;
input x13069;
input x4701;
input x12902;
input x13698;
input x13567;
input x13038;
input x4392;
input x4861;
input x4496;
input x4821;
input x192485;
input x13004;
input x12780;
input x13994;
input x4778;
input x4635;
input x13330;
input x4323;
input x12969;
input x13560;
input x13031;
input x13750;
input x12922;
input x13252;
input x4576;
input x13018;
input x13047;
input x13494;
input x13208;
input x13174;
input x13433;
input x13594;
input x13440;
input x13126;
input x13403;
input x4805;
input x13193;
input x13474;
input x13341;
input x13423;
input x13612;
input x13843;
input x13100;
input x13663;
input x12843;
input x13234;
input x13633;
input x4764;
input x12810;
input x12991;
input x13011;
input x13541;
input x13025;
input x13396;
input x4707;
input x13291;
input x13644;
input x13447;
input x13654;
input x13093;
input x4964;
input x13414;
input x4840;
input x13145;
input x13263;
input x12929;
input x13733;
input x13853;
input x4812;
input x13547;
input x13576;
input x13921;
input x12915;
input x13553;
input x4771;
input x12962;
input x13514;
input x4733;
input x13605;
input x13271;
input x13863;
input x4347;
input x4919;
input x13742;
input x192486;
input x13534;
input x13833;
input x13501;
input x14005;
input x13722;
input x13761;
input x13508;
input x13684;
input x13705;
input x4538;
input x13527;
input x13969;
input x13884;
input x13797;
input x4796;
input x13586;
input x4367;
input x13950;
input x4831;
input x13984;
input x12940;
input x4570;
input x12980;
input x13385;
input x13482;
input x13619;
input x13464;
input x4869;
input x4514;
input x13115;
input x13772;
input x4448;
input x13488;
input x12768;
input x4503;
input x4902;
input x12955;
input x4788;
input x4693;
input x13374;
input x192484;
input x4607;
input x13086;
input x13826;
input x13815;
input x4757;
input x13077;
input x13457;
input x4561;
input x13163;
input x13870;
input x4254;
input x4667;

// Start POs
output x757;
output x749;
output x291;
output x508;
output x971;
output x2633;
output x729;
output x4227;
output x4234;
output x451;
output x1244;
output x815;
output x3122;
output x1087;
output x3996;
output x1032;
output x912;
output x4059;
output x1024;
output x3954;
output x3524;
output x2693;
output x468;
output x378;
output x1215;
output x225;
output x364;
output x3816;
output x852;
output x594;
output x1721;
output x712;
output x2981;
output x1745;
output x879;
output x1062;
output x352;
output x3372;
output x420;
output x1575;
output x4214;
output x4023;
output x827;
output x753;
output x764;
output x697;
output x521;
output x3028;
output x9;
output x4192;
output x3803;
output x3762;
output x170;
output x186;
output x3861;
output x240;
output x845;
output x725;
output x4154;
output x926;
output x4049;
output x132;
output x2594;
output x1152;
output x871;
output x3258;
output x338;
output x3968;
output x2805;
output x863;
output x434;
output x1885;
output x3561;
output x963;
output x4082;
output x52;
output x20;
output x4115;
output x2068;
output x1039;
output x1778;
output x3925;
output x2542;
output x1340;
output x808;
output x0;
output x2308;
output x1977;
output x3418;
output x3604;
output x27;
output x1855;
output x2494;
output x2006;
output x4143;
output x2100;
output x4104;
output x2856;
output x890;
output x1804;
output x2451;
output x3904;
output x3847;
output x3712;
output x608;
output x1829;
output x1174;
output x1532;
output x1383;
output x3485;
output x76;
output x771;
output x831;
output x4070;
output x683;
output x820;
output x1639;
output x1690;
output x2746;
output x306;
output x2908;
output x2400;
output x778;
output x3938;
output x999;
output x3830;
output x3685;
output x3874;
output x480;
output x956;
output x105;
output x1597;
output x2169;
output x801;
output x3451;
output x2355;
output x933;
output x735;
output x4093;
output x649;
output x1912;
output x641;
output x919;
output x661;
output x653;
output x2230;
output x3156;
output x1070;
output x1130;
output x2261;
output x552;
output x677;
output x494;
output x905;
output x3327;
output x1195;
output x785;
output x1305;
output x2948;
output x43;
output x719;
output x668;
output x838;
output x4132;
output x4011;
output x742;
output x154;
output x1016;
output x690;
output x703;
output x4036;
output x563;
output x2041;
output x886;
output x1010;
output x34;
output x394;
output x1281;
output x4166;
output x3207;
output x2133;
output x3079;
output x898;
output x1500;
output x258;
output x324;
output x3288;
output x789;
output x275;
output x1935;
output x1467;
output x3891;
output x208;
output x406;
output x577;
output x1107;
output x1667;
output x1428;
output x794;
output x626;
output x2195;
output x4204;
output x856;
output x4179;
output x3651;
output x3983;
output x534;

// Start wires
wire net_15987;
wire net_8631;
wire net_4065;
wire net_11968;
wire net_4854;
wire net_2418;
wire net_16075;
wire net_7279;
wire net_11788;
wire net_4598;
wire net_12833;
wire net_1897;
wire net_980;
wire net_5499;
wire net_9803;
wire net_12029;
wire net_7081;
wire net_10629;
wire net_11370;
wire net_5515;
wire net_3996;
wire net_18920;
wire net_17083;
wire net_15044;
wire net_6241;
wire net_7298;
wire net_4382;
wire net_13988;
wire net_13226;
wire net_12501;
wire x4861;
wire net_8105;
wire net_4306;
wire net_264;
wire net_12959;
wire net_11178;
wire net_18857;
wire net_3904;
wire net_17256;
wire net_8914;
wire net_17057;
wire net_11757;
wire net_9072;
wire net_2769;
wire net_3707;
wire net_14405;
wire net_2082;
wire net_5035;
wire net_4832;
wire net_4464;
wire net_8577;
wire net_16142;
wire net_17675;
wire net_15913;
wire net_18014;
wire net_703;
wire net_5330;
wire net_193;
wire net_11377;
wire net_9989;
wire net_12447;
wire net_14381;
wire net_6773;
wire net_5273;
wire net_12413;
wire net_16843;
wire net_2942;
wire net_18119;
wire net_13993;
wire net_18314;
wire net_17574;
wire net_13916;
wire net_4442;
wire net_3134;
wire net_13458;
wire net_5523;
wire net_1720;
wire net_14164;
wire net_16825;
wire net_13885;
wire net_8191;
wire net_15098;
wire net_6104;
wire net_2060;
wire net_2051;
wire net_6087;
wire net_4535;
wire net_16807;
wire net_6426;
wire net_593;
wire net_5563;
wire net_10156;
wire net_18422;
wire net_16544;
wire net_6238;
wire net_17216;
wire net_2765;
wire net_15665;
wire net_15085;
wire net_8341;
wire net_18353;
wire net_11044;
wire net_18683;
wire net_16383;
wire net_9597;
wire net_10343;
wire net_15449;
wire net_10320;
wire net_1198;
wire net_3975;
wire net_2862;
wire net_8100;
wire net_2457;
wire net_18237;
wire net_8260;
wire net_5533;
wire net_1516;
wire net_6782;
wire net_6473;
wire net_18777;
wire net_17317;
wire net_1083;
wire net_3423;
wire net_964;
wire net_2913;
wire net_17245;
wire net_16018;
wire net_18257;
wire net_13729;
wire net_6402;
wire net_11003;
wire net_2268;
wire net_17930;
wire net_14352;
wire net_17384;
wire net_17044;
wire net_2846;
wire net_13331;
wire net_11685;
wire net_9479;
wire net_4369;
wire net_18283;
wire net_16364;
wire x12768;
wire net_6401;
wire net_10007;
wire net_4929;
wire net_3959;
wire net_4309;
wire net_8873;
wire net_12393;
wire net_11226;
wire net_6573;
wire net_1140;
wire net_18060;
wire net_2764;
wire net_1464;
wire net_16423;
wire net_11985;
wire net_4973;
wire net_3196;
wire net_14740;
wire net_5962;
wire net_515;
wire net_10620;
wire net_6806;
wire x749;
wire net_5121;
wire net_223;
wire net_15725;
wire net_7146;
wire net_2077;
wire net_15028;
wire net_7496;
wire net_16933;
wire net_2745;
wire net_16856;
wire net_13973;
wire net_5084;
wire net_3965;
wire net_13827;
wire net_15008;
wire net_6706;
wire net_7212;
wire net_572;
wire net_5289;
wire net_10955;
wire net_9614;
wire net_7850;
wire net_1662;
wire net_10396;
wire net_14615;
wire net_1079;
wire net_10148;
wire net_6760;
wire net_5198;
wire net_14318;
wire net_3235;
wire net_4938;
wire net_7099;
wire net_13261;
wire net_2391;
wire net_2802;
wire net_7965;
wire net_4614;
wire net_2906;
wire net_456;
wire net_18332;
wire net_11299;
wire net_7238;
wire net_16750;
wire net_8533;
wire net_3428;
wire net_15781;
wire net_14528;
wire net_493;
wire net_16378;
wire net_6374;
wire net_6080;
wire net_14306;
wire x1778;
wire net_6506;
wire net_987;
wire net_15963;
wire net_6167;
wire net_3620;
wire net_7781;
wire net_13824;
wire net_8475;
wire net_3271;
wire net_13183;
wire net_11197;
wire net_10675;
wire net_13098;
wire net_12568;
wire net_12276;
wire net_12418;
wire net_18816;
wire net_721;
wire net_9033;
wire net_7779;
wire net_8164;
wire net_15590;
wire net_12127;
wire net_13634;
wire net_1018;
wire net_11085;
wire net_11701;
wire net_13289;
wire net_18519;
wire net_6591;
wire net_823;
wire net_9067;
wire net_9269;
wire net_7271;
wire net_4788;
wire net_11774;
wire net_9541;
wire net_7892;
wire net_11028;
wire net_17367;
wire net_5428;
wire net_1191;
wire net_13688;
wire net_16311;
wire net_2255;
wire net_4754;
wire net_17485;
wire net_17596;
wire net_8970;
wire net_16236;
wire net_7471;
wire net_12918;
wire net_16257;
wire net_1019;
wire net_1616;
wire net_17389;
wire net_6180;
wire x653;
wire net_10348;
wire net_16064;
wire net_16625;
wire net_15902;
wire net_9415;
wire net_14181;
wire net_4342;
wire x905;
wire net_12863;
wire net_2969;
wire net_7518;
wire net_12522;
wire net_12351;
wire net_5490;
wire net_12960;
wire net_18734;
wire net_13167;
wire net_15078;
wire net_11406;
wire net_8886;
wire net_2985;
wire net_11551;
wire net_537;
wire net_18750;
wire net_12943;
wire net_11310;
wire net_10893;
wire net_12477;
wire net_13446;
wire net_5501;
wire net_18880;
wire net_12294;
wire net_3252;
wire net_17130;
wire net_18753;
wire net_16184;
wire net_5790;
wire net_5891;
wire net_513;
wire net_12020;
wire net_7950;
wire net_1576;
wire net_1421;
wire net_14282;
wire net_12462;
wire net_17742;
wire net_8737;
wire net_2736;
wire net_1280;
wire net_459;
wire net_12616;
wire net_9239;
wire net_6590;
wire net_18510;
wire net_3412;
wire net_2113;
wire net_13305;
wire net_9397;
wire net_4793;
wire net_4760;
wire net_3915;
wire net_12737;
wire net_14424;
wire net_18938;
wire net_5606;
wire net_8063;
wire net_8353;
wire net_5150;
wire net_9212;
wire net_12713;
wire net_8176;
wire net_11493;
wire net_7709;
wire net_12672;
wire net_18275;
wire net_1659;
wire net_589;
wire net_18329;
wire net_1814;
wire net_17851;
wire net_11610;
wire net_5981;
wire net_16703;
wire net_10186;
wire net_7319;
wire net_8698;
wire net_724;
wire net_9826;
wire net_9123;
wire net_8058;
wire net_2384;
wire net_16784;
wire net_16229;
wire net_7760;
wire net_5889;
wire net_2480;
wire net_9943;
wire net_12181;
wire net_9868;
wire net_874;
wire net_13706;
wire net_15909;
wire net_15264;
wire net_11399;
wire net_4277;
wire net_7907;
wire net_12107;
wire net_3674;
wire net_7555;
wire net_6187;
wire net_4966;
wire net_17749;
wire net_15522;
wire net_14973;
wire net_5244;
wire net_10178;
wire net_11182;
wire net_12857;
wire net_436;
wire net_18713;
wire net_2837;
wire net_7963;
wire net_7181;
wire net_5641;
wire net_11157;
wire net_2824;
wire net_1777;
wire net_12983;
wire net_8263;
wire net_18602;
wire net_15706;
wire net_13647;
wire net_12325;
wire net_7246;
wire net_12153;
wire net_12134;
wire net_5556;
wire net_17534;
wire net_1702;
wire net_4403;
wire net_7974;
wire net_6358;
wire net_16728;
wire net_1838;
wire net_11365;
wire net_10857;
wire net_358;
wire net_1973;
wire net_8748;
wire net_2934;
wire net_11427;
wire net_18026;
wire net_1285;
wire net_10364;
wire net_5912;
wire net_3112;
wire net_15320;
wire net_1175;
wire net_13207;
wire net_13118;
wire x4514;
wire net_9453;
wire net_18361;
wire net_15970;
wire net_9934;
wire net_5722;
wire net_9312;
wire net_9191;
wire net_2922;
wire net_1742;
wire net_11884;
wire net_18003;
wire net_7641;
wire net_17427;
wire x3288;
wire net_11823;
wire net_6890;
wire net_8011;
wire net_17988;
wire net_15368;
wire net_13734;
wire net_3370;
wire net_7025;
wire net_13040;
wire x757;
wire net_15830;
wire net_9497;
wire net_3947;
wire net_3441;
wire net_18213;
wire net_4947;
wire net_16915;
wire net_4015;
wire net_3662;
wire net_12730;
wire net_16586;
wire net_8729;
wire net_9187;
wire net_13441;
wire net_16688;
wire net_6349;
wire net_16451;
wire net_16086;
wire net_10756;
wire net_17879;
wire net_18549;
wire net_3539;
wire net_2031;
wire net_1560;
wire net_4414;
wire net_12451;
wire net_4409;
wire net_17831;
wire net_12160;
wire net_10453;
wire net_6754;
wire net_17870;
wire net_13690;
wire net_8538;
wire net_9684;
wire net_8715;
wire net_14227;
wire net_13111;
wire net_7724;
wire net_6489;
wire net_1545;
wire net_4662;
wire net_18627;
wire net_8204;
wire net_10798;
wire net_18254;
wire net_13838;
wire net_2332;
wire net_12491;
wire net_2715;
wire net_1941;
wire net_14915;
wire net_13074;
wire net_13968;
wire net_14276;
wire net_3899;
wire net_17052;
wire net_1319;
wire net_8757;
wire net_3080;
wire net_11075;
wire net_15091;
wire net_1582;
wire net_4016;
wire net_6028;
wire net_13747;
wire net_2333;
wire net_6544;
wire net_6464;
wire net_17210;
wire net_1368;
wire net_1248;
wire net_2238;
wire net_845;
wire net_10745;
wire net_8003;
wire net_10973;
wire net_9081;
wire net_695;
wire net_18987;
wire net_7692;
wire net_14086;
wire net_2671;
wire net_6787;
wire net_6569;
wire net_12761;
wire net_18542;
wire net_5896;
wire net_12788;
wire net_15169;
wire net_12610;
wire net_14605;
wire net_2198;
wire net_9043;
wire net_16341;
wire net_5250;
wire net_6435;
wire net_6661;
wire net_2940;
wire net_8672;
wire net_16346;
wire net_5583;
wire net_2095;
wire net_4681;
wire net_6955;
wire net_5231;
wire net_9726;
wire net_2314;
wire net_9905;
wire net_5454;
wire net_2613;
wire net_18958;
wire net_15311;
wire net_9995;
wire net_9010;
wire net_8849;
wire net_11479;
wire net_231;
wire net_10197;
wire net_16122;
wire net_17519;
wire net_3024;
wire x34;
wire net_18860;
wire net_4691;
wire net_18520;
wire net_17445;
wire net_12381;
wire net_17110;
wire net_4223;
wire net_11321;
wire net_2297;
wire net_13052;
wire net_9439;
wire net_3325;
wire net_6171;
wire net_582;
wire net_12485;
wire net_16671;
wire net_15331;
wire net_17187;
wire net_7419;
wire net_2341;
wire net_661;
wire net_3360;
wire net_13537;
wire net_15648;
wire net_11854;
wire net_17289;
wire net_9086;
wire net_18461;
wire net_10006;
wire net_9460;
wire net_17165;
wire net_18639;
wire net_210;
wire net_916;
wire net_3395;
wire net_11641;
wire net_4335;
wire net_851;
wire net_9924;
wire net_14865;
wire net_13247;
wire net_2426;
wire net_18196;
wire net_7405;
wire net_12237;
wire net_3310;
wire net_671;
wire net_8817;
wire net_8846;
wire net_14425;
wire net_12431;
wire net_6830;
wire net_6965;
wire net_8734;
wire net_18436;
wire net_16545;
wire net_12978;
wire net_9054;
wire net_17999;
wire net_15473;
wire net_307;
wire net_13938;
wire net_3547;
wire net_14497;
wire net_3543;
wire net_11470;
wire net_15298;
wire net_5104;
wire net_15248;
wire net_14774;
wire net_6069;
wire net_17935;
wire net_2656;
wire net_6326;
wire net_3922;
wire net_3212;
wire net_6530;
wire net_9632;
wire net_1764;
wire net_17684;
wire net_14067;
wire net_3513;
wire net_9968;
wire net_13290;
wire net_4042;
wire net_9691;
wire net_3335;
wire net_5377;
wire net_3682;
wire net_6456;
wire net_18198;
wire net_12245;
wire net_5655;
wire net_18168;
wire net_16839;
wire net_7856;
wire net_2667;
wire net_12818;
wire net_17238;
wire net_5431;
wire net_8443;
wire net_480;
wire net_7662;
wire net_4507;
wire net_4986;
wire net_2897;
wire net_18611;
wire net_5810;
wire x13553;
wire net_836;
wire net_13817;
wire net_18382;
wire net_2161;
wire net_18551;
wire net_12075;
wire net_10671;
wire net_6568;
wire net_8408;
wire net_6059;
wire net_370;
wire net_16470;
wire net_16026;
wire net_13429;
wire net_6443;
wire net_1169;
wire net_13416;
wire net_7057;
wire net_7013;
wire net_13677;
wire net_9238;
wire net_7389;
wire net_2206;
wire net_11206;
wire net_1392;
wire net_14575;
wire net_6121;
wire net_311;
wire net_2479;
wire net_10132;
wire net_15453;
wire net_11119;
wire net_4469;
wire net_11452;
wire net_17726;
wire net_14598;
wire net_16280;
wire net_12527;
wire x13772;
wire net_17899;
wire net_9986;
wire net_13210;
wire net_2520;
wire net_10166;
wire net_10768;
wire net_10704;
wire net_6676;
wire net_2197;
wire net_15943;
wire net_10521;
wire net_5399;
wire net_10220;
wire net_12089;
wire net_9473;
wire net_14658;
wire net_2905;
wire net_10372;
wire net_200;
wire net_4435;
wire net_16489;
wire net_16032;
wire net_8612;
wire net_5220;
wire net_16463;
wire net_5995;
wire net_16208;
wire net_14706;
wire net_1853;
wire net_9741;
wire net_10119;
wire net_10240;
wire net_2170;
wire net_6851;
wire net_15304;
wire net_15026;
wire net_2678;
wire net_17605;
wire net_11036;
wire net_8346;
wire net_9119;
wire net_16965;
wire net_10256;
wire net_8906;
wire net_6698;
wire net_18228;
wire net_11267;
wire net_18301;
wire net_10381;
wire net_15609;
wire net_7717;
wire net_6988;
wire net_6281;
wire net_6209;
wire net_2864;
wire net_1998;
wire net_9341;
wire net_13621;
wire net_11656;
wire net_2795;
wire net_13587;
wire net_5540;
wire net_16214;
wire net_16166;
wire net_1918;
wire net_12790;
wire net_18421;
wire net_15388;
wire net_5870;
wire net_7894;
wire net_3236;
wire net_17964;
wire net_5837;
wire net_3201;
wire net_11812;
wire net_11169;
wire net_8147;
wire net_8096;
wire net_5613;
wire net_17510;
wire net_9560;
wire net_8966;
wire net_7163;
wire net_17889;
wire net_8024;
wire net_6897;
wire net_12912;
wire net_5300;
wire net_12359;
wire net_8926;
wire net_18677;
wire x0;
wire net_5803;
wire net_5410;
wire net_14838;
wire net_3650;
wire net_2465;
wire net_15544;
wire net_5078;
wire net_5447;
wire net_12043;
wire net_15230;
wire net_14465;
wire net_8485;
wire net_10388;
wire net_7462;
wire net_9900;
wire net_6023;
wire net_13862;
wire net_898;
wire x13447;
wire net_14855;
wire net_6136;
wire net_10416;
wire net_16288;
wire net_15548;
wire net_13023;
wire net_8364;
wire net_7229;
wire net_7045;
wire net_8640;
wire net_1376;
wire net_5005;
wire net_13409;
wire net_8810;
wire net_6885;
wire net_6701;
wire net_18792;
wire net_1980;
wire net_13793;
wire net_9303;
wire net_1302;
wire net_244;
wire net_7341;
wire x3451;
wire net_8687;
wire net_2395;
wire net_6012;
wire net_5347;
wire net_5439;
wire net_4002;
wire net_1989;
wire net_18642;
wire net_2855;
wire net_1795;
wire net_13310;
wire net_9247;
wire net_18878;
wire net_12186;
wire net_17597;
wire net_1539;
wire net_9626;
wire net_16538;
wire net_17193;
wire net_4261;
wire net_18871;
wire net_10123;
wire net_3490;
wire net_3035;
wire net_7646;
wire net_14417;
wire net_15191;
wire net_11483;
wire net_13434;
wire net_16100;
wire net_6359;
wire net_12082;
wire net_11131;
wire net_7430;
wire net_7437;
wire net_1469;
wire net_15749;
wire net_11626;
wire net_18927;
wire net_4081;
wire net_15694;
wire net_2436;
wire net_18427;
wire net_16811;
wire net_16403;
wire net_16454;
wire net_10793;
wire net_14176;
wire net_11878;
wire net_621;
wire net_10018;
wire net_5153;
wire net_13316;
wire net_10375;
wire net_12586;
wire net_18246;
wire net_7729;
wire net_5598;
wire net_12591;
wire net_11276;
wire net_3985;
wire net_14492;
wire net_18648;
wire net_14801;
wire net_12390;
wire net_9792;
wire x3954;
wire net_18770;
wire net_9552;
wire net_10229;
wire net_9689;
wire net_18101;
wire net_12663;
wire net_13032;
wire net_999;
wire net_15783;
wire net_8549;
wire net_10888;
wire net_8838;
wire net_13924;
wire net_9752;
wire net_4994;
wire net_3588;
wire net_9151;
wire net_1480;
wire net_18912;
wire net_14759;
wire net_15839;
wire net_7700;
wire net_4952;
wire net_377;
wire net_8836;
wire net_288;
wire net_16640;
wire net_2649;
wire net_1459;
wire net_12252;
wire net_7290;
wire net_5265;
wire net_11650;
wire x13193;
wire net_7749;
wire net_3741;
wire net_13257;
wire net_4470;
wire net_9168;
wire net_540;
wire net_2642;
wire net_6650;
wire net_891;
wire net_12899;
wire net_9388;
wire net_5224;
wire net_3065;
wire net_5821;
wire net_4167;
wire net_15011;
wire net_7796;
wire net_6746;
wire net_4711;
wire net_10236;
wire net_5868;
wire net_18059;
wire net_10358;
wire net_18336;
wire net_16437;
wire net_4802;
wire net_16635;
wire net_618;
wire net_18786;
wire net_9075;
wire net_3688;
wire net_5759;
wire net_12001;
wire net_12399;
wire net_8256;
wire net_6970;
wire net_14907;
wire net_14255;
wire net_5945;
wire net_6148;
wire net_754;
wire net_10785;
wire net_7193;
wire net_921;
wire net_9113;
wire net_7989;
wire net_17569;
wire net_11581;
wire net_4957;
wire net_14900;
wire net_3308;
wire net_12607;
wire net_10274;
wire net_16772;
wire net_2192;
wire net_1533;
wire net_16440;
wire net_16336;
wire net_8565;
wire net_7999;
wire net_7681;
wire net_9138;
wire net_15525;
wire net_11158;
wire net_9884;
wire net_3502;
wire net_14014;
wire net_4827;
wire net_654;
wire net_17248;
wire net_330;
wire net_3506;
wire net_16953;
wire net_8082;
wire net_14538;
wire net_9116;
wire net_570;
wire net_444;
wire net_525;
wire net_3829;
wire net_3646;
wire net_1210;
wire net_1067;
wire net_15575;
wire net_6624;
wire net_5058;
wire net_18746;
wire net_16882;
wire net_14920;
wire net_5998;
wire net_7820;
wire net_16971;
wire net_14681;
wire net_16569;
wire x4166;
wire net_6200;
wire net_6259;
wire net_15206;
wire net_3933;
wire net_18584;
wire net_11629;
wire net_16300;
wire net_9325;
wire net_4820;
wire x3651;
wire net_13486;
wire net_10055;
wire net_7577;
wire net_16579;
wire net_15828;
wire net_9409;
wire net_9404;
wire net_1178;
wire net_9722;
wire net_5573;
wire net_17372;
wire net_7098;
wire net_3825;
wire net_11142;
wire net_6218;
wire net_17177;
wire net_16097;
wire net_12380;
wire net_340;
wire net_6039;
wire net_16057;
wire net_15885;
wire net_15435;
wire net_2634;
wire net_434;
wire net_6915;
wire net_8434;
wire net_7024;
wire net_6936;
wire net_14200;
wire net_1797;
wire net_9443;
wire net_11086;
wire net_14732;
wire net_4906;
wire net_4524;
wire net_339;
wire net_7686;
wire net_17848;
wire net_13105;
wire net_3468;
wire net_10443;
wire net_11775;
wire net_18918;
wire net_12753;
wire net_2710;
wire net_15722;
wire net_2660;
wire net_14486;
wire net_8624;
wire net_10083;
wire net_8087;
wire net_5389;
wire net_3671;
wire net_8236;
wire net_8651;
wire net_3691;
wire net_17562;
wire net_678;
wire net_15771;
wire net_16503;
wire net_11631;
wire net_8979;
wire net_928;
wire net_15251;
wire net_5459;
wire net_13363;
wire net_208;
wire net_9225;
wire net_7878;
wire net_8215;
wire net_2744;
wire net_2377;
wire net_415;
wire net_3251;
wire net_2786;
wire net_347;
wire net_14784;
wire net_13526;
wire net_11059;
wire net_3794;
wire x820;
wire net_12664;
wire net_15997;
wire net_7306;
wire net_16551;
wire net_1335;
wire net_18874;
wire net_15716;
wire net_15519;
wire net_12210;
wire net_5477;
wire net_18154;
wire net_16932;
wire net_2212;
wire net_5453;
wire net_11535;
wire net_7730;
wire net_16725;
wire x1912;
wire net_16499;
wire net_3571;
wire net_4642;
wire net_610;
wire net_8130;
wire net_16889;
wire net_7870;
wire net_15187;
wire net_2344;
wire net_10588;
wire net_1323;
wire net_14130;
wire net_1506;
wire net_10470;
wire net_17836;
wire net_13386;
wire net_6496;
wire net_13193;
wire net_539;
wire net_16617;
wire net_13068;
wire net_692;
wire net_16094;
wire net_18971;
wire net_4568;
wire net_10807;
wire net_17551;
wire net_4377;
wire net_16660;
wire net_15130;
wire net_14261;
wire net_7704;
wire net_13125;
wire net_15104;
wire net_10311;
wire net_1400;
wire net_885;
wire net_9202;
wire net_11698;
wire net_14320;
wire net_9918;
wire net_18276;
wire net_10770;
wire net_6822;
wire net_11607;
wire net_6594;
wire net_3517;
wire net_761;
wire net_496;
wire net_11396;
wire net_1554;
wire net_7101;
wire net_16779;
wire net_10638;
wire net_4370;
wire net_18980;
wire net_4979;
wire net_14613;
wire net_12578;
wire net_2249;
wire net_16106;
wire net_5686;
wire net_15129;
wire net_739;
wire x5001;
wire net_8760;
wire net_17529;
wire net_17472;
wire net_826;
wire net_15069;
wire net_1738;
wire net_10384;
wire net_10504;
wire net_14887;
wire net_16178;
wire net_11644;
wire net_6716;
wire net_2624;
wire net_11761;
wire net_343;
wire net_17038;
wire net_7313;
wire net_9672;
wire net_8456;
wire net_5236;
wire net_4424;
wire net_7541;
wire net_9615;
wire net_7451;
wire net_2487;
wire net_7803;
wire net_8227;
wire net_17649;
wire net_13132;
wire net_15674;
wire net_2975;
wire net_17201;
wire net_4625;
wire net_5257;
wire net_8220;
wire net_2779;
wire net_14187;
wire net_11552;
wire net_17494;
wire net_16225;
wire net_6392;
wire net_18990;
wire net_15158;
wire net_9346;
wire net_11352;
wire net_8169;
wire net_1490;
wire net_9274;
wire net_4282;
wire net_15216;
wire net_17066;
wire net_11806;
wire net_12774;
wire net_18923;
wire net_17926;
wire net_15565;
wire net_14765;
wire net_14342;
wire net_5742;
wire net_4356;
wire net_685;
wire net_8466;
wire net_18808;
wire net_16307;
wire net_12349;
wire net_17711;
wire net_11843;
wire net_4052;
wire net_8513;
wire net_18224;
wire net_8681;
wire net_15953;
wire x1639;
wire net_16897;
wire net_17049;
wire net_13469;
wire net_10652;
wire net_7160;
wire net_17633;
wire net_12876;
wire net_4686;
wire net_1946;
wire net_2733;
wire net_17204;
wire net_14280;
wire net_18697;
wire net_6764;
wire net_13252;
wire net_6769;
wire net_3612;
wire net_11634;
wire net_1605;
wire net_12795;
wire net_18726;
wire net_18702;
wire net_5118;
wire net_747;
wire net_15597;
wire net_2305;
wire net_1653;
wire net_14125;
wire net_5842;
wire net_9817;
wire net_7377;
wire net_16023;
wire net_2258;
wire net_11168;
wire net_12510;
wire net_14327;
wire net_17397;
wire net_6500;
wire net_17276;
wire net_2367;
wire net_15977;
wire net_14697;
wire net_4573;
wire net_4127;
wire net_16900;
wire net_2810;
wire net_13546;
wire net_1053;
wire net_11292;
wire net_1004;
wire net_4921;
wire net_17939;
wire net_11716;
wire net_11359;
wire net_3232;
wire net_13356;
wire net_4498;
wire net_3228;
wire net_2282;
wire net_10029;
wire net_1546;
wire net_11367;
wire net_8542;
wire net_15695;
wire net_6042;
wire net_13654;
wire net_18849;
wire net_16390;
wire net_1046;
wire net_19016;
wire net_11502;
wire net_10332;
wire net_4960;
wire net_1213;
wire net_2265;
wire net_8118;
wire net_16948;
wire net_10163;
wire net_16479;
wire net_5795;
wire net_12812;
wire net_769;
wire net_1780;
wire net_13668;
wire net_16132;
wire net_1025;
wire net_3758;
wire net_15062;
wire net_13157;
wire net_10403;
wire net_7502;
wire net_15807;
wire net_1089;
wire net_12169;
wire net_16359;
wire net_11998;
wire net_16386;
wire net_4528;
wire net_6233;
wire net_5625;
wire net_16695;
wire net_4141;
wire net_18292;
wire net_14094;
wire net_12535;
wire net_10669;
wire net_5146;
wire net_16713;
wire net_8701;
wire net_5326;
wire x4764;
wire net_12921;
wire net_17923;
wire net_4394;
wire net_18082;
wire net_15421;
wire net_5953;
wire net_12442;
wire net_11047;
wire net_12702;
wire net_9433;
wire net_10816;
wire net_14124;
wire net_13248;
wire net_3626;
wire net_15924;
wire net_12095;
wire net_5779;
wire net_14798;
wire net_6417;
wire net_4726;
wire net_15475;
wire net_14377;
wire net_13086;
wire net_9588;
wire net_18033;
wire net_17220;
wire net_14572;
wire net_5344;
wire net_7492;
wire net_12468;
wire net_5364;
wire net_18945;
wire net_8743;
wire net_6388;
wire net_13478;
wire net_740;
wire net_4072;
wire net_11090;
wire net_5825;
wire net_3183;
wire net_17863;
wire net_3908;
wire net_4837;
wire net_730;
wire net_4150;
wire net_8049;
wire net_7094;
wire net_5405;
wire net_11931;
wire net_2105;
wire net_16371;
wire net_7226;
wire net_1127;
wire net_6381;
wire net_17226;
wire net_9458;
wire net_11243;
wire net_6420;
wire net_13831;
wire net_18176;
wire net_7465;
wire net_9297;
wire net_15732;
wire net_4143;
wire net_12900;
wire net_18768;
wire net_8679;
wire net_7285;
wire x13797;
wire net_5140;
wire net_3123;
wire net_2955;
wire net_771;
wire net_2301;
wire net_2978;
wire net_15033;
wire net_5185;
wire net_13139;
wire net_3950;
wire net_1062;
wire net_14395;
wire net_4936;
wire net_3293;
wire net_4120;
wire net_9246;
wire net_7733;
wire net_16263;
wire net_14987;
wire net_6050;
wire net_13214;
wire net_5188;
wire net_4590;
wire net_18343;
wire net_18096;
wire net_6116;
wire net_16512;
wire net_1411;
wire net_12549;
wire net_505;
wire net_4088;
wire net_16862;
wire net_10471;
wire net_3723;
wire net_14724;
wire net_10493;
wire net_10426;
wire net_7152;
wire net_6527;
wire net_992;
wire net_7485;
wire net_15933;
wire net_9781;
wire net_6727;
wire net_782;
wire net_10527;
wire net_13576;
wire net_11106;
wire net_18347;
wire net_6291;
wire net_4186;
wire net_13328;
wire net_4738;
wire net_3314;
wire net_7422;
wire net_2971;
wire net_5776;
wire net_17102;
wire net_13322;
wire net_10339;
wire net_8072;
wire net_8244;
wire net_2836;
wire net_10615;
wire net_5689;
wire net_7429;
wire net_1805;
wire net_4667;
wire net_11536;
wire net_10660;
wire net_3635;
wire net_17838;
wire net_13559;
wire net_7120;
wire net_1110;
wire net_17423;
wire net_15356;
wire net_442;
wire net_14999;
wire net_13789;
wire net_16594;
wire net_7202;
wire net_3087;
wire net_17402;
wire net_14627;
wire net_13900;
wire net_1821;
wire x4082;
wire net_11675;
wire net_7480;
wire net_3865;
wire net_1588;
wire net_9029;
wire net_4037;
wire net_3937;
wire net_1495;
wire net_17080;
wire net_18800;
wire net_2992;
wire net_12974;
wire net_17227;
wire net_16329;
wire net_3522;
wire x3847;
wire net_668;
wire net_7601;
wire net_18142;
wire net_15758;
wire net_3079;
wire net_14203;
wire net_17733;
wire net_8040;
wire net_5814;
wire net_12707;
wire net_1070;
wire net_8878;
wire net_1225;
wire net_812;
wire x999;
wire net_14993;
wire net_13805;
wire net_18830;
wire net_6314;
wire net_6972;
wire net_1107;
wire net_16563;
wire net_15850;
wire net_11053;
wire net_18581;
wire net_15621;
wire net_3384;
wire net_1203;
wire net_13347;
wire net_15055;
wire net_9011;
wire net_12402;
wire net_12176;
wire net_10867;
wire net_10715;
wire net_5321;
wire net_11434;
wire net_12789;
wire net_17440;
wire net_17652;
wire net_5884;
wire net_863;
wire net_7131;
wire net_6468;
wire net_3164;
wire net_16527;
wire net_16998;
wire net_14058;
wire net_13150;
wire net_904;
wire net_15580;
wire net_12850;
wire net_14226;
wire net_13552;
wire net_16244;
wire net_6777;
wire net_12286;
wire net_6633;
wire net_8126;
wire net_6092;
wire net_16813;
wire net_6559;
wire net_15553;
wire net_11360;
wire net_9183;
wire net_15688;
wire net_4845;
wire net_1160;
wire net_18630;
wire net_15917;
wire net_159;
wire net_11147;
wire net_9379;
wire net_3268;
wire net_18939;
wire net_5863;
wire net_11615;
wire net_9523;
wire net_10181;
wire net_9354;
wire net_14834;
wire net_2875;
wire net_12952;
wire net_10213;
wire x4743;
wire net_324;
wire net_6848;
wire net_11724;
wire net_10284;
wire net_10074;
wire net_13397;
wire net_5480;
wire net_14675;
wire net_10309;
wire net_18761;
wire net_16354;
wire net_7257;
wire net_17776;
wire net_13047;
wire net_9706;
wire x4023;
wire net_14248;
wire net_14103;
wire net_17616;
wire net_12647;
wire net_10964;
wire net_5046;
wire net_3066;
wire net_6270;
wire net_15385;
wire net_6275;
wire net_17805;
wire net_4181;
wire net_376;
wire net_17909;
wire net_2133;
wire net_17703;
wire net_13643;
wire net_16978;
wire net_4817;
wire net_13374;
wire net_2515;
wire net_19020;
wire net_3173;
wire net_8038;
wire net_3738;
wire net_17393;
wire net_7994;
wire net_15529;
wire net_5298;
wire net_5119;
wire net_422;
wire net_4290;
wire net_18048;
wire net_14739;
wire net_1345;
wire net_1450;
wire net_561;
wire net_12694;
wire net_4899;
wire net_5955;
wire net_8501;
wire net_4299;
wire net_2290;
wire net_12741;
wire net_2851;
wire net_17140;
wire net_8427;
wire net_14640;
wire net_14019;
wire net_3772;
wire net_7901;
wire net_4868;
wire net_2698;
wire net_6552;
wire net_18653;
wire net_8453;
wire net_3450;
wire net_14412;
wire net_14813;
wire net_3528;
wire net_8559;
wire net_18005;
wire net_8956;
wire x3830;
wire net_350;
wire net_4270;
wire net_8332;
wire net_13178;
wire net_7606;
wire net_13275;
wire net_18075;
wire net_3117;
wire net_16753;
wire net_14245;
wire net_11816;
wire net_3482;
wire net_6648;
wire net_7375;
wire net_15712;
wire net_3369;
wire net_9020;
wire net_1101;
wire net_994;
wire net_12828;
wire net_12268;
wire net_18919;
wire net_6685;
wire net_11837;
wire net_4166;
wire net_4608;
wire net_15122;
wire net_3340;
wire net_4545;
wire net_3844;
wire net_1849;
wire net_10045;
wire net_5486;
wire net_16647;
wire net_13516;
wire net_14994;
wire net_14637;
wire net_11122;
wire net_1108;
wire net_8583;
wire net_9756;
wire net_1878;
wire net_16598;
wire net_16820;
wire net_16231;
wire net_17314;
wire net_13070;
wire net_16678;
wire net_9255;
wire net_16435;
wire net_11446;
wire net_3890;
wire net_5975;
wire net_7528;
wire net_4025;
wire net_16112;
wire net_9194;
wire net_15459;
wire net_7078;
wire x6501;
wire net_7008;
wire net_11957;
wire net_3882;
wire net_557;
wire net_3043;
wire net_15288;
wire net_7860;
wire net_6611;
wire net_13891;
wire net_11386;
wire net_12316;
wire net_1991;
wire net_1611;
wire net_18201;
wire net_14046;
wire net_1431;
wire x879;
wire net_1714;
wire net_18135;
wire net_13014;
wire net_11970;
wire net_16945;
wire net_18827;
wire net_8868;
wire net_240;
wire net_15115;
wire net_15872;
wire net_18147;
wire net_17261;
wire net_17588;
wire net_295;
wire net_8411;
wire net_18558;
wire net_13425;
wire net_9241;
wire net_5935;
wire net_17326;
wire net_13490;
wire net_7753;
wire net_15236;
wire net_14879;
wire net_12115;
wire net_7720;
wire net_16462;
wire net_11239;
wire net_12619;
wire net_6691;
wire net_12967;
wire net_278;
wire net_18208;
wire net_6864;
wire net_19029;
wire net_9063;
wire net_4874;
wire net_10090;
wire net_16794;
wire net_13309;
wire net_17952;
wire net_2443;
wire net_10736;
wire net_1307;
wire net_4514;
wire net_15857;
wire net_17499;
wire net_15753;
wire net_6940;
wire net_5591;
wire net_4810;
wire net_15413;
wire net_4418;
wire net_17959;
wire net_5385;
wire net_14145;
wire net_6099;
wire net_9786;
wire net_12679;
wire net_7630;
wire net_13854;
wire x13705;
wire net_13712;
wire net_3776;
wire net_17954;
wire net_1252;
wire net_9173;
wire net_7739;
wire net_9095;
wire net_7784;
wire net_16700;
wire net_10731;
wire net_507;
wire net_10097;
wire net_8981;
wire net_1902;
wire net_17115;
wire net_7111;
wire net_2600;
wire net_5734;
wire net_3563;
wire net_12224;
wire net_8726;
wire net_6585;
wire net_9565;
wire net_11936;
wire net_4491;
wire net_11543;
wire net_8282;
wire net_7538;
wire net_16737;
wire net_1962;
wire net_291;
wire net_9502;
wire net_7351;
wire net_1964;
wire net_857;
wire net_867;
wire net_5964;
wire net_15618;
wire net_396;
wire x4179;
wire net_14845;
wire net_10602;
wire net_17468;
wire net_8851;
wire net_10535;
wire net_1541;
wire net_14966;
wire net_14216;
wire net_9748;
wire net_15683;
wire net_5177;
wire net_271;
wire net_3329;
wire net_10067;
wire net_6111;
wire net_12208;
wire net_14693;
wire net_3611;
wire net_2064;
wire net_15274;
wire net_5333;
wire net_1925;
wire x594;
wire net_1909;
wire x4392;
wire net_16664;
wire net_1410;
wire net_365;
wire net_13412;
wire net_18043;
wire net_3344;
wire net_12060;
wire net_8374;
wire net_10729;
wire net_4413;
wire net_13849;
wire net_8719;
wire net_4313;
wire net_16483;
wire net_16830;
wire net_11000;
wire net_16448;
wire net_8313;
wire net_16630;
wire net_9339;
wire net_7128;
wire net_7915;
wire x13208;
wire net_13723;
wire net_13730;
wire net_4892;
wire net_803;
wire net_10884;
wire x434;
wire net_14713;
wire net_14111;
wire net_7764;
wire net_6375;
wire net_17501;
wire net_1476;
wire net_1293;
wire net_14939;
wire net_11098;
wire net_2883;
wire net_8665;
wire net_11742;
wire net_2681;
wire x4707;
wire net_12159;
wire net_9629;
wire net_18181;
wire net_17791;
wire net_5136;
wire net_18598;
wire net_4855;
wire net_14668;
wire x13644;
wire net_1266;
wire net_1452;
wire net_2773;
wire net_17995;
wire net_909;
wire net_4529;
wire net_4898;
wire net_152;
wire net_11575;
wire net_3105;
wire net_2138;
wire net_16153;
wire net_258;
wire net_11192;
wire net_10761;
wire net_16196;
wire net_12935;
wire net_12054;
wire net_19033;
wire net_19017;
wire net_13983;
wire net_5083;
wire net_2446;
wire net_18576;
wire net_7171;
wire net_11999;
wire net_15644;
wire net_7605;
wire net_585;
wire net_7611;
wire net_17754;
wire net_7809;
wire net_14823;
wire net_11913;
wire net_11347;
wire net_12061;
wire net_10593;
wire net_14514;
wire net_10293;
wire net_12632;
wire net_788;
wire net_9090;
wire net_214;
wire net_8113;
wire net_13028;
wire net_8144;
wire net_3578;
wire net_12455;
wire net_13903;
wire net_8804;
wire net_6310;
wire net_5097;
wire net_7329;
wire net_18409;
wire net_4259;
wire net_2565;
wire net_17890;
wire net_8018;
wire net_13229;
wire net_6783;
wire net_5908;
wire net_2118;
wire net_463;
wire net_15281;
wire net_17946;
wire net_9487;
wire net_197;
wire net_18867;
wire net_2560;
wire net_9331;
wire net_5017;
wire net_3709;
wire net_13085;
wire net_12803;
wire net_7588;
wire net_11468;
wire net_5352;
wire net_2595;
wire net_1383;
wire net_7302;
wire net_2751;
wire net_9663;
wire net_9165;
wire net_18462;
wire net_4446;
wire net_14160;
wire net_10484;
wire net_6269;
wire net_6176;
wire net_14170;
wire net_13672;
wire net_11116;
wire net_13497;
wire net_1683;
wire net_17178;
wire net_17027;
wire net_12515;
wire net_978;
wire net_15510;
wire net_1313;
wire net_7618;
wire net_3331;
wire net_15855;
wire net_16891;
wire x2693;
wire net_11994;
wire net_13286;
wire net_5712;
wire net_14446;
wire net_10877;
wire net_8383;
wire net_9954;
wire net_6360;
wire net_17351;
wire net_17298;
wire net_1789;
wire net_14035;
wire net_13142;
wire net_13940;
wire net_3219;
wire net_7520;
wire net_4587;
wire net_18286;
wire net_2576;
wire net_2352;
wire net_1038;
wire net_6931;
wire net_4241;
wire net_9920;
wire net_8168;
wire net_5710;
wire net_5369;
wire net_3763;
wire net_15445;
wire net_6333;
wire net_11338;
wire net_14662;
wire net_7697;
wire net_2277;
wire net_17162;
wire net_6078;
wire net_975;
wire net_5421;
wire net_15538;
wire net_4650;
wire net_15805;
wire net_13061;
wire net_15735;
wire net_6160;
wire net_5874;
wire net_18489;
wire net_2006;
wire net_13570;
wire net_1331;
wire net_18474;
wire net_12307;
wire net_15071;
wire net_5826;
wire net_18908;
wire net_13912;
wire net_18065;
wire net_16071;
wire net_8604;
wire net_2728;
wire net_17070;
wire net_18109;
wire net_4636;
wire net_6264;
wire net_17991;
wire net_13619;
wire net_12847;
wire net_11514;
wire net_10026;
wire net_16550;
wire net_9262;
wire net_18456;
wire net_14752;
wire x2169;
wire net_4092;
wire net_17406;
wire net_12300;
wire net_8595;
wire net_11760;
wire net_10751;
wire net_15361;
wire net_4486;
wire net_9427;
wire net_18054;
wire net_9131;
wire net_15905;
wire net_17197;
wire net_10983;
wire net_7262;
wire net_387;
wire net_15327;
wire net_3275;
wire net_7447;
wire net_6297;
wire net_18524;
wire net_17660;
wire net_10828;
wire net_5291;
wire net_1893;
wire net_16509;
wire net_15355;
wire net_1932;
wire net_9639;
wire net_8896;
wire net_11620;
wire net_8268;
wire net_3836;
wire net_15777;
wire net_14554;
wire net_1957;
wire net_10102;
wire net_13743;
wire net_13231;
wire net_9368;
wire net_15377;
wire net_7581;
wire net_2572;
wire net_2414;
wire net_19003;
wire net_1846;
wire x1935;
wire net_13381;
wire net_5667;
wire net_11222;
wire net_9662;
wire net_7888;
wire net_12475;
wire net_11066;
wire net_13984;
wire x534;
wire net_4254;
wire net_13760;
wire net_3815;
wire net_3555;
wire net_17810;
wire net_18538;
wire net_5739;
wire net_2371;
wire net_6794;
wire net_14077;
wire net_13368;
wire net_11014;
wire net_16622;
wire net_8396;
wire net_12546;
wire net_9640;
wire net_7843;
wire net_7392;
wire net_3982;
wire net_1388;
wire net_4709;
wire net_14409;
wire net_14959;
wire x13038;
wire net_9858;
wire net_3391;
wire net_15018;
wire net_2730;
wire net_6835;
wire net_13553;
wire net_4655;
wire net_1624;
wire net_6618;
wire net_12332;
wire net_1638;
wire net_7455;
wire net_3875;
wire net_12146;
wire net_9319;
wire net_14436;
wire net_10135;
wire net_5268;
wire net_11389;
wire net_14980;
wire net_6335;
wire net_2153;
wire net_17692;
wire net_1939;
wire net_9582;
wire net_8781;
wire net_3098;
wire net_7242;
wire net_14190;
wire net_6288;
wire net_4673;
wire net_5762;
wire net_9061;
wire net_10249;
wire net_16852;
wire net_7828;
wire net_162;
wire net_15751;
wire net_14952;
wire net_8301;
wire net_7776;
wire net_653;
wire net_14301;
wire net_13160;
wire net_16909;
wire net_5066;
wire net_13919;
wire net_14718;
wire net_11735;
wire net_12030;
wire x2006;
wire net_3145;
wire net_9558;
wire net_15879;
wire net_13694;
wire net_3694;
wire net_16001;
wire net_18661;
wire net_14880;
wire net_10262;
wire net_11592;
wire net_3855;
wire net_236;
wire net_12324;
wire net_9286;
wire net_552;
wire net_10823;
wire net_8206;
wire net_1787;
wire net_17897;
wire net_3551;
wire net_6654;
wire net_7440;
wire net_14791;
wire net_13390;
wire net_9518;
wire net_7067;
wire net_17300;
wire net_16980;
wire net_15143;
wire net_16910;
wire net_8329;
wire net_14402;
wire net_3416;
wire net_7198;
wire net_18686;
wire net_5166;
wire net_17609;
wire net_15992;
wire net_14595;
wire net_4886;
wire net_9878;
wire net_17479;
wire net_15655;
wire net_10914;
wire net_14070;
wire net_12039;
wire net_8522;
wire net_6659;
wire net_12192;
wire net_6877;
wire net_711;
wire net_17882;
wire net_15635;
wire net_18952;
wire net_17309;
wire net_8618;
wire net_4700;
wire net_846;
wire net_17152;
wire net_3017;
wire net_11864;
wire net_4677;
wire net_16880;
wire net_8033;
wire net_16515;
wire net_10996;
wire net_10038;
wire net_5768;
wire net_18021;
wire net_2607;
wire net_7799;
wire net_15210;
wire net_7957;
wire net_10971;
wire net_14755;
wire net_8769;
wire net_13870;
wire net_5023;
wire net_2168;
wire net_18072;
wire net_17091;
wire net_1885;
wire net_1030;
wire net_14357;
wire net_10406;
wire net_6929;
wire net_16272;
wire net_10682;
wire net_15498;
wire net_11498;
wire net_10031;
wire net_4773;
wire net_4201;
wire net_4273;
wire net_1969;
wire net_7991;
wire net_15514;
wire net_12306;
wire net_8009;
wire net_7064;
wire net_17007;
wire net_933;
wire net_12532;
wire net_12036;
wire net_10860;
wire net_3377;
wire net_373;
wire net_16573;
wire net_16357;
wire x1024;
wire net_452;
wire net_16046;
wire net_3683;
wire net_1483;
wire net_8067;
wire net_3031;
wire net_17707;
wire net_2645;
wire net_10433;
wire net_5356;
wire net_14386;
wire net_8078;
wire net_7674;
wire net_7386;
wire net_6684;
wire net_4278;
wire net_2674;
wire net_16847;
wire net_13801;
wire net_10193;
wire net_8934;
wire net_7059;
wire net_14428;
wire net_1671;
wire net_4764;
wire net_665;
wire net_1746;
wire net_2222;
wire net_2825;
wire net_17343;
wire net_7209;
wire net_18478;
wire net_3670;
wire net_14647;
wire net_5940;
wire net_5985;
wire net_7925;
wire net_16565;
wire net_6606;
wire net_10182;
wire net_10376;
wire net_4861;
wire net_11666;
wire net_1706;
wire net_16691;
wire net_3574;
wire net_18796;
wire net_5994;
wire net_10852;
wire net_2921;
wire net_3289;
wire net_8829;
wire net_10225;
wire net_3114;
wire net_3415;
wire net_10019;
wire net_744;
wire net_16430;
wire net_8276;
wire net_15620;
wire net_18430;
wire net_17530;
wire net_7985;
wire net_4136;
wire net_2011;
wire net_15023;
wire net_777;
wire net_4806;
wire net_13203;
wire net_7185;
wire net_3157;
wire net_7532;
wire net_490;
wire net_18297;
wire net_17746;
wire net_14805;
wire net_11497;
wire net_12677;
wire net_18782;
wire net_12130;
wire net_13930;
wire net_6009;
wire net_3462;
wire net_5670;
wire net_4439;
wire net_5602;
wire net_7638;
wire net_2841;
wire net_10106;
wire net_11889;
wire net_7255;
wire net_5813;
wire net_1977;
wire net_2938;
wire net_14009;
wire net_14568;
wire net_1171;
wire net_10691;
wire net_9680;
wire net_248;
wire net_3594;
wire net_17989;
wire net_6548;
wire net_5341;
wire net_16995;
wire net_16562;
wire net_14064;
wire net_13583;
wire net_15268;
wire net_18616;
wire net_18580;
wire net_1767;
wire net_4010;
wire net_7333;
wire net_11827;
wire net_1640;
wire net_12956;
wire net_13788;
wire net_2724;
wire net_11916;
wire net_12090;
wire net_15762;
wire net_1741;
wire net_16708;
wire net_10141;
wire net_16163;
wire net_4227;
wire net_7550;
wire net_959;
wire net_5381;
wire net_11476;
wire net_7911;
wire net_3051;
wire net_2345;
wire net_6981;
wire net_16643;
wire net_6460;
wire net_6660;
wire net_2164;
wire net_11079;
wire net_5659;
wire net_11797;
wire net_3751;
wire x13808;
wire net_5311;
wire net_4564;
wire net_2338;
wire net_15685;
wire net_2616;
wire net_8200;
wire net_282;
wire net_1596;
wire net_17039;
wire net_10804;
wire net_4296;
wire x753;
wire net_11857;
wire net_10908;
wire net_11693;
wire net_2370;
wire net_2047;
wire net_8320;
wire net_9647;
wire net_12733;
wire net_2693;
wire net_13115;
wire net_11212;
wire net_16711;
wire net_12765;
wire net_12185;
wire net_9621;
wire net_907;
wire net_18909;
wire net_14473;
wire net_3076;
wire net_16103;
wire net_2719;
wire net_6343;
wire net_9688;
wire net_16126;
wire net_641;
wire net_2798;
wire net_5071;
wire net_10977;
wire net_3869;
wire net_14335;
wire net_1152;
wire net_1226;
wire net_14212;
wire net_10525;
wire net_5315;
wire net_15533;
wire net_14976;
wire net_10257;
wire net_3805;
wire net_15865;
wire net_16764;
wire net_3942;
wire net_15823;
wire net_15352;
wire net_7836;
wire net_13199;
wire net_1818;
wire net_12783;
wire net_11850;
wire net_13335;
wire net_8646;
wire net_9371;
wire net_17013;
wire net_1523;
wire net_1656;
wire net_17095;
wire net_6522;
wire net_16315;
wire net_17558;
wire net_15179;
wire net_691;
wire net_6951;
wire net_5551;
wire net_3178;
wire net_2701;
wire net_17356;
wire net_10422;
wire net_1863;
wire net_15108;
wire net_10774;
wire net_8399;
wire net_2519;
wire net_471;
wire net_18210;
wire net_18000;
wire net_1055;
wire net_3894;
wire net_878;
wire net_518;
wire net_11136;
wire net_10172;
wire net_14523;
wire net_13533;
wire net_929;
wire net_18853;
wire net_17045;
wire x4132;
wire net_2523;
wire net_11779;
wire net_4210;
wire net_3954;
wire net_12939;
wire net_11811;
wire net_5726;
wire net_1565;
wire net_5262;
wire net_14487;
wire net_169;
wire net_17738;
wire net_15347;
wire net_9948;
wire net_16869;
wire net_12986;
wire net_2234;
wire net_16318;
wire net_12120;
wire net_17000;
wire net_15629;
wire net_17727;
wire net_6828;
wire net_10481;
wire net_967;
wire net_13056;
wire net_4420;
wire net_8007;
wire net_13861;
wire net_4318;
wire net_12358;
wire net_11475;
wire net_4910;
wire net_17172;
wire net_1645;
wire net_2962;
wire net_16428;
wire net_4365;
wire net_176;
wire net_12410;
wire net_15036;
wire net_614;
wire net_17570;
wire net_12505;
wire net_8293;
wire net_3194;
wire net_3572;
wire net_5537;
wire net_4740;
wire net_8338;
wire net_1192;
wire net_10697;
wire net_6857;
wire net_14368;
wire net_4542;
wire net_11753;
wire net_11705;
wire net_15093;
wire net_8730;
wire net_4061;
wire net_12201;
wire net_3156;
wire net_12109;
wire net_2482;
wire net_13043;
wire net_7275;
wire net_707;
wire net_6534;
wire net_5039;
wire net_11174;
wire net_6867;
wire net_18038;
wire net_18175;
wire net_4850;
wire net_13828;
wire net_4531;
wire net_14778;
wire net_575;
wire net_5833;
wire net_18184;
wire net_4715;
wire net_7169;
wire net_3697;
wire net_18993;
wire net_11374;
wire net_14810;
wire net_12582;
wire net_6193;
wire net_16188;
wire net_15962;
wire net_6431;
wire net_3618;
wire net_9156;
wire net_7562;
wire net_15893;
wire net_14012;
wire net_10842;
wire net_16829;
wire net_5512;
wire net_765;
wire net_1342;
wire net_2633;
wire net_1666;
wire net_4193;
wire net_15661;
wire net_8573;
wire net_8253;
wire net_17249;
wire net_2099;
wire net_15390;
wire net_5745;
wire net_6750;
wire net_5182;
wire net_7612;
wire net_18757;
wire net_13454;
wire net_18088;
wire net_16659;
wire net_9809;
wire net_10302;
wire net_17679;
wire net_16308;
wire net_16137;
wire net_8195;
wire net_5850;
wire net_5646;
wire net_2021;
wire net_11248;
wire net_1068;
wire net_186;
wire net_2495;
wire net_15229;
wire net_12823;
wire net_6672;
wire net_16803;
wire x3938;
wire net_1050;
wire net_17670;
wire net_2760;
wire net_5914;
wire net_4751;
wire net_15910;
wire net_2271;
wire net_5327;
wire net_16036;
wire net_14083;
wire net_18902;
wire net_12164;
wire net_6125;
wire net_7143;
wire net_16014;
wire net_7983;
wire net_10324;
wire net_3130;
wire net_8572;
wire net_15157;
wire net_16478;
wire net_17340;
wire net_5704;
wire x12980;
wire net_4289;
wire net_9775;
wire x742;
wire net_9510;
wire net_13806;
wire net_4712;
wire net_11340;
wire net_260;
wire net_2947;
wire net_15729;
wire net_12552;
wire net_11784;
wire net_3137;
wire net_8649;
wire net_12423;
wire net_1597;
wire net_16911;
wire net_7946;
wire net_8785;
wire net_7593;
wire net_3988;
wire x1107;
wire net_17056;
wire net_2761;
wire net_6396;
wire net_3788;
wire net_15605;
wire net_4355;
wire net_16007;
wire net_10623;
wire net_1503;
wire net_3961;
wire net_8430;
wire net_4639;
wire net_8628;
wire net_11089;
wire net_5494;
wire net_9299;
wire net_17885;
wire net_11928;
wire net_9574;
wire net_12638;
wire net_9606;
wire net_12362;
wire net_11409;
wire net_6595;
wire net_13663;
wire net_11653;
wire net_13866;
wire net_17362;
wire net_5443;
wire net_5211;
wire net_4731;
wire net_2989;
wire net_497;
wire net_6720;
wire net_12494;
wire net_7658;
wire net_15291;
wire net_8160;
wire net_1414;
wire net_4153;
wire net_11307;
wire net_10927;
wire net_9864;
wire net_300;
wire net_2652;
wire net_5526;
wire net_10149;
wire net_1233;
wire net_2720;
wire net_6351;
wire net_15058;
wire net_12917;
wire net_1834;
wire net_6027;
wire net_4925;
wire net_17285;
wire net_13213;
wire net_15258;
wire net_13024;
wire net_13313;
wire net_15690;
wire net_11355;
wire net_5474;
wire net_14363;
wire net_9745;
wire net_8984;
wire net_12565;
wire net_15888;
wire net_13405;
wire net_10203;
wire net_11946;
wire net_13603;
wire net_5194;
wire net_12025;
wire net_3150;
wire net_9596;
wire net_15967;
wire net_3979;
wire net_8822;
wire net_15927;
wire net_12712;
wire net_839;
wire net_13542;
wire net_11778;
wire net_7095;
wire net_18754;
wire net_4660;
wire net_13013;
wire net_17719;
wire net_18504;
wire net_11294;
wire net_7805;
wire net_11313;
wire net_954;
wire net_18415;
wire net_13094;
wire x192486;
wire net_4565;
wire net_9051;
wire net_9037;
wire net_15048;
wire net_8796;
wire net_11271;
wire net_8962;
wire net_10897;
wire net_16957;
wire net_16412;
wire net_10152;
wire x4538;
wire net_15671;
wire net_16253;
wire net_13359;
wire net_13265;
wire net_14456;
wire net_9545;
wire net_10411;
wire net_18730;
wire net_12445;
wire net_11989;
wire net_4790;
wire net_12048;
wire net_17383;
wire net_5363;
wire net_7529;
wire net_8888;
wire net_6665;
wire net_16921;
wire net_4900;
wire net_9807;
wire net_13222;
wire net_6502;
wire net_14888;
wire net_14783;
wire net_7305;
wire net_6163;
wire net_3011;
wire net_17577;
wire net_13079;
wire net_10643;
wire net_18229;
wire net_13187;
wire net_10021;
wire net_12946;
wire net_6817;
wire net_6000;
wire net_9079;
wire net_8863;
wire net_14859;
wire net_11930;
wire net_13628;
wire net_12466;
wire net_9536;
wire net_17592;
wire net_12887;
wire net_3010;
wire net_881;
wire net_12657;
wire net_17877;
wire net_10544;
wire net_2805;
wire net_1397;
wire net_14619;
wire net_14231;
wire net_15182;
wire net_4474;
wire net_18373;
wire net_14623;
wire net_17566;
wire net_16290;
wire net_1954;
wire net_13036;
wire net_7615;
wire net_17272;
wire net_14294;
wire net_14924;
wire net_2041;
wire net_17933;
wire net_13090;
wire net_16628;
wire net_11830;
wire net_10354;
wire net_7937;
wire net_18056;
wire net_7930;
wire net_7196;
wire net_16613;
wire net_12197;
wire net_14143;
wire net_2423;
wire net_7535;
wire net_6723;
wire net_13875;
wire net_12379;
wire net_11283;
wire net_895;
wire net_10781;
wire net_6412;
wire net_18475;
wire net_14469;
wire net_11603;
wire net_5990;
wire net_14358;
wire net_15202;
wire net_12006;
wire net_8240;
wire net_7048;
wire net_9715;
wire net_7767;
wire net_17683;
wire net_8831;
wire net_12394;
wire net_10683;
wire net_1255;
wire net_12603;
wire net_1250;
wire net_8247;
wire net_13928;
wire net_16395;
wire net_15176;
wire net_16937;
wire net_207;
wire net_3643;
wire net_18743;
wire net_19045;
wire net_15149;
wire net_16775;
wire net_13639;
wire net_17782;
wire net_12102;
wire net_13382;
wire net_11874;
wire net_1689;
wire net_10345;
wire net_10271;
wire net_6186;
wire net_17783;
wire net_15466;
wire net_8569;
wire net_5698;
wire net_274;
wire net_13987;
wire net_1075;
wire net_9387;
wire net_13360;
wire net_6204;
wire net_930;
wire net_2387;
wire net_12599;
wire net_9316;
wire net_8358;
wire net_4723;
wire net_2267;
wire net_7323;
wire net_4769;
wire net_18217;
wire net_16740;
wire net_13590;
wire x956;
wire net_10016;
wire net_4888;
wire net_9539;
wire net_18013;
wire net_14636;
wire net_17528;
wire net_19008;
wire net_3304;
wire net_15382;
wire net_2549;
wire net_11024;
wire net_8654;
wire net_14390;
wire x4367;
wire net_3465;
wire net_18658;
wire net_6217;
wire net_637;
wire net_15787;
wire net_13062;
wire net_2390;
wire net_5436;
wire net_2686;
wire net_5577;
wire net_1509;
wire net_529;
wire net_18493;
wire net_9447;
wire net_3495;
wire net_9887;
wire net_2553;
wire net_17548;
wire net_4881;
wire net_18113;
wire net_8506;
wire net_6477;
wire net_11303;
wire net_16076;
wire net_5228;
wire net_7475;
wire net_15324;
wire net_16305;
wire net_16908;
wire net_9762;
wire net_15579;
wire net_3820;
wire net_3799;
wire net_4175;
wire net_10938;
wire net_2664;
wire net_18403;
wire net_14206;
wire net_11202;
wire net_849;
wire net_14161;
wire net_17563;
wire net_10577;
wire net_7470;
wire net_5294;
wire net_11681;
wire net_14545;
wire net_5751;
wire net_401;
wire net_8165;
wire net_17376;
wire net_10720;
wire net_3798;
wire net_14906;
wire net_2714;
wire net_2183;
wire net_2557;
wire net_14903;
wire net_14265;
wire net_9229;
wire net_11361;
wire x12902;
wire net_758;
wire net_14955;
wire net_13754;
wire net_6874;
wire net_14482;
wire net_10846;
wire net_13563;
wire net_7682;
wire net_5504;
wire net_18233;
wire net_15133;
wire net_4998;
wire net_3255;
wire net_12303;
wire net_9848;
wire net_6564;
wire net_16052;
wire net_15835;
wire net_9797;
wire net_12973;
wire net_10946;
wire net_16098;
wire net_5306;
wire net_9577;
wire net_9938;
wire net_11539;
wire net_16893;
wire net_2917;
wire net_8404;
wire net_15630;
wire net_6711;
wire net_3221;
wire net_16936;
wire net_7708;
wire net_605;
wire net_3411;
wire net_4987;
wire net_10447;
wire net_17291;
wire net_9233;
wire net_9527;
wire net_924;
wire net_8883;
wire net_12255;
wire net_17323;
wire net_5469;
wire net_9205;
wire net_10980;
wire net_16444;
wire net_7829;
wire net_2348;
wire net_489;
wire net_14911;
wire net_17476;
wire net_5457;
wire net_6143;
wire net_4646;
wire net_18774;
wire net_2748;
wire net_9991;
wire net_18150;
wire net_11561;
wire net_9611;
wire net_9135;
wire net_8060;
wire net_251;
wire net_15772;
wire net_840;
wire net_9206;
wire x4093;
wire net_10632;
wire net_8086;
wire net_17845;
wire net_6933;
wire net_15429;
wire net_5789;
wire net_13281;
wire net_12928;
wire net_11229;
wire net_9914;
wire net_411;
wire net_2137;
wire net_11689;
wire net_15075;
wire net_12220;
wire net_11256;
wire net_12688;
wire net_7874;
wire net_7293;
wire net_8975;
wire net_1862;
wire net_13889;
wire net_10052;
wire net_2317;
wire net_6248;
wire net_16118;
wire net_8135;
wire net_16885;
wire x13385;
wire net_10584;
wire net_6035;
wire net_6492;
wire net_3583;
wire net_8183;
wire net_19030;
wire net_10536;
wire net_8219;
wire net_15802;
wire net_2373;
wire net_11694;
wire net_14109;
wire net_17310;
wire net_16332;
wire net_10943;
wire net_7746;
wire net_9282;
wire net_15137;
wire net_1609;
wire net_402;
wire net_7847;
wire net_4047;
wire net_3448;
wire net_7108;
wire net_3248;
wire net_12450;
wire net_2274;
wire net_11597;
wire net_12681;
wire net_17602;
wire net_11488;
wire net_13859;
wire net_10950;
wire net_18842;
wire net_12345;
wire x2633;
wire net_2359;
wire net_16835;
wire net_15038;
wire net_16701;
wire net_13101;
wire net_12574;
wire net_15432;
wire net_11585;
wire net_16473;
wire net_10127;
wire net_4102;
wire net_6908;
wire net_1430;
wire net_9964;
wire net_6892;
wire net_2478;
wire net_6429;
wire net_2563;
wire net_18040;
wire net_12435;
wire net_9484;
wire net_9243;
wire net_8051;
wire net_5679;
wire net_16729;
wire net_3408;
wire net_4870;
wire net_630;
wire net_12514;
wire net_2202;
wire net_2490;
wire net_8841;
wire net_14861;
wire net_4428;
wire net_1791;
wire net_4339;
wire net_1471;
wire net_9975;
wire net_8997;
wire net_7667;
wire net_3608;
wire net_18079;
wire net_17088;
wire net_16602;
wire net_14892;
wire net_912;
wire net_17034;
wire net_13562;
wire net_7018;
wire net_4517;
wire net_15315;
wire net_3841;
wire net_1928;
wire net_1328;
wire net_9871;
wire net_16458;
wire net_2859;
wire net_3848;
wire net_2884;
wire net_5372;
wire net_4942;
wire net_13616;
wire net_3205;
wire net_1094;
wire net_3487;
wire net_2749;
wire net_855;
wire net_674;
wire net_18935;
wire net_11032;
wire net_9506;
wire net_303;
wire net_10041;
wire net_15821;
wire net_18647;
wire net_9982;
wire net_2475;
wire net_9925;
wire net_18328;
wire net_2937;
wire net_7792;
wire net_7657;
wire net_7400;
wire net_6191;
wire net_17168;
wire net_14744;
wire net_12249;
wire net_16746;
wire net_12993;
wire net_7865;
wire net_4743;
wire net_13767;
wire net_17960;
wire net_9478;
wire net_2439;
wire net_13297;
wire net_11048;
wire net_172;
wire net_4341;
wire net_13460;
wire net_15300;
wire net_4048;
wire net_17234;
wire net_16962;
wire net_10749;
wire net_4570;
wire net_17832;
wire net_16284;
wire net_10244;
wire net_18449;
wire net_6689;
wire x13684;
wire net_12233;
wire net_13934;
wire net_7034;
wire net_6446;
wire net_8029;
wire net_11939;
wire net_9050;
wire net_6198;
wire net_3733;
wire net_3881;
wire net_12263;
wire net_8598;
wire net_11944;
wire net_10519;
wire net_14136;
wire net_15481;
wire net_8091;
wire net_8057;
wire net_6258;
wire net_8361;
wire net_1758;
wire net_13840;
wire net_8813;
wire net_18571;
wire net_16549;
wire net_14868;
wire net_11802;
wire net_1769;
wire net_9115;
wire net_6694;
wire net_15504;
wire net_1567;
wire net_17940;
wire net_8020;
wire net_6322;
wire net_12087;
wire net_15286;
wire net_11186;
wire net_8152;
wire net_18193;
wire net_9520;
wire net_14930;
wire net_476;
wire net_2783;
wire net_17513;
wire net_14461;
wire net_6055;
wire net_7079;
wire net_382;
wire net_11412;
wire net_11259;
wire net_5301;
wire net_583;
wire net_7041;
wire net_16987;
wire net_15947;
wire net_9408;
wire net_17996;
wire net_14173;
wire net_16734;
wire net_17967;
wire net_13055;
wire net_9695;
wire net_4719;
wire net_17071;
wire net_10379;
wire net_17827;
wire net_15234;
wire net_9005;
wire net_4460;
wire net_220;
wire net_1465;
wire net_11153;
wire net_13599;
wire net_4982;
wire net_16407;
wire net_543;
wire net_625;
wire net_3760;
wire net_17469;
wire net_16944;
wire net_11411;
wire net_10708;
wire net_17796;
wire net_15543;
wire net_17506;
wire net_11637;
wire net_14509;
wire net_13790;
wire net_4331;
wire net_2909;
wire net_4953;
wire net_15464;
wire net_9607;
wire net_4697;
wire net_5638;
wire net_7899;
wire net_15594;
wire net_12157;
wire net_10562;
wire net_1694;
wire net_12844;
wire x12810;
wire net_4991;
wire net_910;
wire net_15940;
wire net_12356;
wire net_15332;
wire net_18514;
wire net_5394;
wire net_7944;
wire x3418;
wire net_2412;
wire net_16247;
wire x4104;
wire net_12070;
wire net_4265;
wire net_18717;
wire net_14563;
wire net_4158;
wire net_13442;
wire net_17078;
wire net_13527;
wire net_315;
wire net_1375;
wire net_18411;
wire net_4006;
wire net_16969;
wire net_8212;
wire net_1351;
wire net_17455;
wire net_18673;
wire net_1535;
wire net_16859;
wire net_2400;
wire net_5543;
wire net_18261;
wire x13547;
wire net_8661;
wire net_10959;
wire net_2034;
wire net_15189;
wire net_14963;
wire net_8921;
wire net_1808;
wire net_3256;
wire net_13122;
wire net_18164;
wire net_15003;
wire net_14916;
wire net_13438;
wire net_10567;
wire net_3322;
wire net_2533;
wire net_10267;
wire net_1913;
wire net_12297;
wire net_16024;
wire net_13243;
wire net_11526;
wire net_7830;
wire net_16413;
wire net_9673;
wire net_9016;
wire net_7642;
wire net_11904;
wire net_9732;
wire net_9264;
wire net_15244;
wire net_6615;
wire net_12279;
wire net_7409;
wire net_7671;
wire net_1760;
wire net_7714;
wire net_3926;
wire net_4849;
wire net_5758;
wire net_3403;
wire net_10002;
wire net_6977;
wire net_10718;
wire net_3093;
wire net_7935;
wire net_12820;
wire net_6886;
wire net_647;
wire net_3247;
wire net_15745;
wire net_17975;
wire net_18962;
wire net_6452;
wire net_8684;
wire net_2464;
wire net_12272;
wire net_9492;
wire net_3839;
wire net_6513;
wire net_17722;
wire net_17349;
wire net_2732;
wire net_13483;
wire net_11809;
wire net_8368;
wire net_7345;
wire net_1096;
wire net_795;
wire net_8153;
wire net_18425;
wire net_11403;
wire net_1406;
wire net_9093;
wire net_15754;
wire net_18965;
wire net_8490;
wire net_18986;
wire net_10463;
wire net_1434;
wire net_6996;
wire net_3668;
wire net_14728;
wire net_6096;
wire x4851;
wire net_9823;
wire net_10012;
wire net_5130;
wire net_11870;
wire net_5617;
wire net_4946;
wire net_774;
wire net_15101;
wire net_18804;
wire net_10071;
wire net_6958;
wire net_8892;
wire net_13235;
wire net_7221;
wire net_501;
wire net_3679;
wire net_4489;
wire net_12344;
wire net_5818;
wire net_6213;
wire net_4692;
wire net_9769;
wire net_6644;
wire net_7481;
wire net_9170;
wire net_13327;
wire net_447;
wire net_9180;
wire net_15126;
wire net_13279;
wire net_5772;
wire net_6318;
wire net_11219;
wire net_14031;
wire net_10755;
wire net_16590;
wire net_13371;
wire net_9703;
wire net_12368;
wire net_8952;
wire net_13944;
wire net_10923;
wire net_7900;
wire net_18563;
wire net_14038;
wire net_4106;
wire net_2951;
wire net_8621;
wire net_3631;
wire net_12854;
wire x2308;
wire net_18707;
wire net_2293;
wire net_16681;
wire net_10105;
wire net_1802;
wire net_15100;
wire net_7694;
wire net_5482;
wire net_10456;
wire net_7637;
wire net_11318;
wire net_18045;
wire net_2755;
wire net_12172;
wire x683;
wire net_13850;
wire net_1678;
wire net_14997;
wire net_6638;
wire net_3366;
wire net_10210;
wire net_15338;
wire net_18628;
wire net_8271;
wire net_7737;
wire net_7206;
wire net_6757;
wire net_17656;
wire net_8511;
wire net_7757;
wire net_11726;
wire net_15442;
wire net_10934;
wire net_3436;
wire net_18069;
wire net_18136;
wire net_14159;
wire net_15500;
wire net_10812;
wire net_8708;
wire net_7725;
wire net_3911;
wire net_17441;
wire net_13913;
wire net_12866;
wire net_5337;
wire net_15557;
wire net_8638;
wire net_17929;
wire net_3365;
wire net_10711;
wire net_18390;
wire net_14372;
wire net_14099;
wire net_12698;
wire net_8587;
wire net_1114;
wire net_10619;
wire net_13431;
wire net_7090;
wire net_3388;
wire net_10664;
wire net_4116;
wire net_3218;
wire net_18386;
wire net_13005;
wire net_4632;
wire net_12283;
wire net_18525;
wire net_8171;
wire net_7266;
wire net_6738;
wire net_18700;
wire net_6690;
wire net_6565;
wire net_18559;
wire net_3811;
wire net_1028;
wire net_14287;
wire net_1529;
wire net_600;
wire net_14021;
wire net_397;
wire net_11126;
wire net_7602;
wire net_5595;
wire net_10968;
wire net_9894;
wire net_12373;
wire net_1384;
wire net_17518;
wire net_17181;
wire net_8712;
wire net_3918;
wire net_9107;
wire net_5280;
wire net_320;
wire net_6844;
wire net_16240;
wire net_4916;
wire net_6902;
wire net_15211;
wire net_9251;
wire net_9103;
wire net_12530;
wire net_7063;
wire net_986;
wire net_1242;
wire x13058;
wire net_15980;
wire net_6556;
wire net_4346;
wire net_1241;
wire net_15571;
wire net_13153;
wire net_11953;
wire net_3690;
wire net_15584;
wire net_7524;
wire net_11833;
wire net_11019;
wire net_13998;
wire net_13197;
wire net_17581;
wire net_3001;
wire net_3121;
wire net_10368;
wire net_4841;
wire net_4621;
wire net_10289;
wire net_10217;
wire net_1634;
wire net_10305;
wire net_6271;
wire net_609;
wire net_12034;
wire net_13343;
wire net_6155;
wire net_3083;
wire net_5693;
wire net_17612;
wire net_9782;
wire net_1221;
wire net_15419;
wire net_7158;
wire net_6911;
wire net_4895;
wire net_9851;
wire net_14943;
wire net_816;
wire net_16005;
wire net_16082;
wire net_9100;
wire net_3264;
wire net_7363;
wire net_2092;
wire net_16872;
wire net_13209;
wire net_7134;
wire net_12745;
wire net_8669;
wire net_18230;
wire net_1217;
wire net_13879;
wire net_7028;
wire net_9719;
wire net_2933;
wire net_8141;
wire net_3381;
wire net_10818;
wire net_16344;
wire net_14156;
wire net_8848;
wire net_18895;
wire net_4118;
wire net_4577;
wire net_17913;
wire net_4970;
wire net_1575;
wire net_17821;
wire net_3279;
wire net_657;
wire net_8495;
wire net_5042;
wire net_1727;
wire net_17644;
wire net_16367;
wire net_329;
wire net_16757;
wire net_5809;
wire net_4600;
wire net_14633;
wire net_12848;
wire net_1924;
wire net_4287;
wire net_1825;
wire net_3168;
wire net_16674;
wire net_10078;
wire net_14714;
wire net_10558;
wire net_962;
wire net_7914;
wire net_8695;
wire net_13731;
wire net_7817;
wire net_596;
wire net_11840;
wire net_1261;
wire net_2120;
wire net_15081;
wire net_4705;
wire net_10430;
wire net_14167;
wire net_7566;
wire net_14735;
wire net_13512;
wire net_18657;
wire net_12893;
wire net_565;
wire net_2569;
wire net_2832;
wire net_4478;
wire net_2149;
wire net_18904;
wire net_13174;
wire net_9736;
wire net_15654;
wire net_10611;
wire net_17304;
wire net_10363;
wire net_16785;
wire net_5062;
wire net_6518;
wire net_4236;
wire net_11618;
wire net_17772;
wire net_18372;
wire net_4813;
wire net_14679;
wire net_10986;
wire net_232;
wire net_16260;
wire net_6538;
wire net_14273;
wire net_18787;
wire net_12778;
wire net_2167;
wire net_2880;
wire net_16350;
wire net_15408;
wire net_7923;
wire net_11062;
wire net_2996;
wire net_6386;
wire net_15147;
wire net_4465;
wire net_532;
wire net_2501;
wire net_3530;
wire net_13179;
wire net_14751;
wire net_14817;
wire net_18516;
wire net_8223;
wire net_889;
wire net_12609;
wire net_1116;
wire x1721;
wire net_13018;
wire net_16879;
wire net_5253;
wire net_17542;
wire net_4373;
wire net_13135;
wire net_9289;
wire net_17498;
wire net_18832;
wire net_11521;
wire net_2814;
wire net_689;
wire net_751;
wire net_16294;
wire net_15172;
wire net_15222;
wire net_14670;
wire net_2363;
wire net_14346;
wire x13174;
wire net_15882;
wire net_3659;
wire net_6578;
wire net_5232;
wire net_13708;
wire net_10512;
wire net_3724;
wire net_13129;
wire net_16556;
wire net_16174;
wire net_4593;
wire net_15615;
wire net_15561;
wire net_1426;
wire net_12649;
wire net_11111;
wire net_9813;
wire net_1407;
wire net_3147;
wire net_4903;
wire net_15343;
wire net_5409;
wire net_12949;
wire net_16043;
wire net_3263;
wire net_10093;
wire net_14610;
wire net_16941;
wire net_14129;
wire net_17137;
wire net_4931;
wire net_16548;
wire net_17715;
wire net_10509;
wire net_7261;
wire net_8613;
wire net_8233;
wire net_6189;
wire net_5114;
wire net_15920;
wire net_4398;
wire net_1042;
wire net_4783;
wire net_4076;
wire net_15703;
wire net_7788;
wire net_17409;
wire net_1000;
wire net_1995;
wire net_17208;
wire net_2545;
wire net_18979;
wire net_5158;
wire net_17751;
wire net_2870;
wire net_14769;
wire net_18358;
wire net_6182;
wire net_4320;
wire net_11847;
wire net_2596;
wire net_10835;
wire net_2970;
wire net_14388;
wire net_12369;
wire net_18117;
wire net_14001;
wire net_9001;
wire net_2584;
wire net_16279;
wire net_14052;
wire net_17764;
wire net_18099;
wire net_18451;
wire net_7546;
wire net_11963;
wire net_952;
wire net_14305;
wire net_4097;
wire net_11743;
wire net_5170;
wire net_3185;
wire net_19025;
wire net_17433;
wire net_13821;
wire net_14290;
wire net_9048;
wire net_3300;
wire net_6438;
wire net_2245;
wire net_7268;
wire net_12963;
wire net_8187;
wire net_7570;
wire net_13773;
wire net_4231;
wire net_383;
wire net_4068;
wire net_14055;
wire net_3140;
wire net_15625;
wire net_6765;
wire net_18500;
wire net_16203;
wire net_427;
wire net_7823;
wire net_1121;
wire net_18123;
wire net_13687;
wire net_7288;
wire net_13897;
wire net_7559;
wire net_18809;
wire net_7381;
wire net_4329;
wire net_16904;
wire net_11094;
wire net_6409;
wire net_2777;
wire net_17464;
wire net_1049;
wire net_13531;
wire net_9440;
wire net_3901;
wire net_17867;
wire net_10674;
wire net_18693;
wire net_14674;
wire net_9364;
wire net_6707;
wire net_8437;
wire net_9278;
wire net_7582;
wire net_6229;
wire net_8608;
wire net_5199;
wire net_12905;
wire net_12388;
wire net_9293;
wire net_18739;
wire net_2591;
wire net_14534;
wire net_10552;
wire net_8985;
wire net_10880;
wire net_17789;
wire net_5189;
wire net_11896;
wire net_5791;
wire net_3968;
wire net_1283;
wire net_16652;
wire net_12875;
wire net_4554;
wire net_18885;
wire net_354;
wire net_14607;
wire net_17067;
wire net_12428;
wire net_15001;
wire net_16267;
wire net_15973;
wire net_18017;
wire net_12099;
wire net_3356;
wire net_11423;
wire net_7175;
wire net_5465;
wire net_12640;
wire net_3886;
wire net_7281;
wire net_1592;
wire net_13650;
wire net_2085;
wire net_4406;
wire net_17416;
wire net_16668;
wire net_12557;
wire net_5621;
wire net_15425;
wire net_8764;
wire net_10297;
wire net_1637;
wire net_3702;
wire net_9374;
wire net_6480;
wire net_6425;
wire net_5971;
wire net_6220;
wire x4070;
wire net_16639;
wire net_8915;
wire net_7629;
wire net_18315;
wire net_11324;
wire net_5854;
wire net_14519;
wire net_4555;
wire net_2070;
wire net_11661;
wire net_16389;
wire net_10605;
wire net_4124;
wire net_16191;
wire net_18934;
wire net_16698;
wire x1597;
wire net_12372;
wire net_3981;
wire net_13659;
wire net_3161;
wire net_6107;
wire net_4303;
wire net_1290;
wire net_12924;
wire net_4147;
wire net_4056;
wire net_17337;
wire net_12589;
wire net_3297;
wire net_14028;
wire net_11766;
wire net_5249;
wire net_13474;
wire net_12205;
wire net_3424;
wire net_18941;
wire net_15371;
wire net_6364;
wire net_10169;
wire net_5087;
wire net_13218;
wire net_11983;
wire net_15397;
wire net_3104;
wire net_5508;
wire net_15066;
wire net_2278;
wire net_3072;
wire net_15409;
wire net_7286;
wire net_1021;
wire net_18680;
wire net_10498;
wire net_5269;
wire net_10488;
wire net_1737;
wire net_9979;
wire net_16375;
wire net_10657;
wire net_6801;
wire net_3607;
wire net_4654;
wire net_8541;
wire net_4917;
wire net_1145;
wire net_8424;
wire net_9306;
wire net_2261;
wire net_9411;
wire net_18949;
wire net_3061;
wire net_7414;
wire net_2958;
wire net_11328;
wire net_14131;
wire net_5918;
wire net_18105;
wire net_10827;
wire net_15869;
wire net_16069;
wire net_6853;
wire net_13961;
wire net_13624;
wire net_6307;
wire net_4192;
wire net_11977;
wire net_14586;
wire net_17330;
wire net_11733;
wire net_11141;
wire net_11568;
wire net_4583;
wire net_18488;
wire net_18222;
wire net_12290;
wire net_4663;
wire net_14330;
wire net_5822;
wire net_4084;
wire net_4500;
wire net_8045;
wire net_15351;
wire net_8591;
wire net_5879;
wire net_14250;
wire net_15812;
wire net_8562;
wire net_2056;
wire net_5716;
wire net_17293;
wire net_7884;
wire net_12217;
wire net_10800;
wire net_9147;
wire net_1628;
wire net_3476;
wire net_15162;
wire net_13957;
wire net_7347;
wire net_4823;
wire net_12519;
wire net_2512;
wire net_12997;
wire net_1936;
wire net_3802;
wire net_14749;
wire net_18219;
wire net_10035;
wire net_14339;
wire net_2708;
wire net_8773;
wire net_8705;
wire net_18996;
wire net_17523;
wire net_10873;
wire net_9958;
wire net_2211;
wire net_18279;
wire net_7425;
wire net_5479;
wire net_16050;
wire net_13001;
wire net_14090;
wire net_8388;
wire net_8777;
wire net_9998;
wire net_1732;
wire net_5926;
wire net_7866;
wire net_6348;
wire net_18485;
wire net_9390;
wire net_12149;
wire net_900;
wire net_7597;
wire net_5528;
wire net_2001;
wire net_1491;
wire net_10879;
wire net_14442;
wire net_8306;
wire net_10918;
wire net_5390;
wire net_18527;
wire net_1034;
wire net_11559;
wire net_16218;
wire net_15634;
wire net_11510;
wire x13984;
wire net_17758;
wire net_17437;
wire net_3439;
wire net_18323;
wire net_13332;
wire net_18159;
wire net_11398;
wire net_1959;
wire net_18212;
wire net_15372;
wire x4902;
wire net_11506;
wire net_12320;
wire net_14884;
wire net_17667;
wire net_460;
wire net_7356;
wire net_6797;
wire net_6074;
wire net_4206;
wire x1428;
wire net_16983;
wire net_15566;
wire net_15365;
wire net_1133;
wire net_15797;
wire net_14788;
wire net_14222;
wire net_6131;
wire net_17062;
wire net_11712;
wire net_10724;
wire net_166;
wire net_14429;
wire net_11027;
wire net_13954;
wire net_5489;
wire net_13164;
wire net_3871;
wire net_18915;
wire net_4455;
wire net_10995;
wire net_8788;
wire net_3352;
wire net_18634;
wire net_7507;
wire net_3832;
wire net_17119;
wire net_5663;
wire net_6017;
wire net_10062;
wire net_17688;
wire net_6925;
wire net_334;
wire net_10930;
wire net_2453;
wire net_3062;
wire net_9586;
wire net_5738;
wire net_12629;
wire net_10952;
wire net_13797;
wire net_16539;
wire net_18364;
wire net_12626;
wire net_14042;
wire net_6790;
wire net_3768;
wire net_2286;
wire net_16716;
wire net_1552;
wire net_13785;
wire net_9380;
wire net_14833;
wire net_14015;
wire net_17556;
wire net_14539;
wire net_5674;
wire net_14532;
wire net_14591;
wire net_7954;
wire x13423;
wire net_3215;
wire net_298;
wire net_1933;
wire net_3717;
wire net_998;
wire net_12620;
wire net_4657;
wire net_2157;
wire net_8945;
wire net_15491;
wire net_10317;
wire net_11154;
wire net_13148;
wire net_12457;
wire net_9328;
wire net_13763;
wire net_14194;
wire net_2405;
wire net_14929;
wire net_835;
wire net_7459;
wire net_15381;
wire net_18592;
wire net_13683;
wire net_9321;
wire net_10466;
wire net_6459;
wire net_17905;
wire net_14795;
wire net_638;
wire net_17916;
wire net_5633;
wire net_18978;
wire net_10028;
wire net_5766;
wire net_11519;
wire net_12801;
wire x4812;
wire net_1783;
wire net_7771;
wire net_1874;
wire net_9554;
wire net_14948;
wire net_14308;
wire net_17251;
wire net_14447;
wire net_3499;
wire net_5206;
wire net_4777;
wire net_17972;
wire net_13192;
wire net_14108;
wire net_12808;
wire net_785;
wire net_9152;
wire net_16490;
wire net_5883;
wire net_4215;
wire net_17920;
wire net_9874;
wire net_6677;
wire net_10902;
wire net_13633;
wire net_10409;
wire net_9657;
wire net_7479;
wire net_3746;
wire net_1349;
wire net_979;
wire net_156;
wire net_13251;
wire net_11820;
wire net_12563;
wire net_2015;
wire net_6658;
wire x4869;
wire net_9676;
wire net_5202;
wire net_4877;
wire net_4170;
wire net_3101;
wire net_12336;
wire net_6268;
wire net_12723;
wire x4788;
wire net_3876;
wire x258;
wire net_16576;
wire net_5982;
wire net_1887;
wire net_13146;
wire net_7444;
wire net_5470;
wire net_14851;
wire net_4033;
wire net_4245;
wire net_11868;
wire net_9514;
wire net_5568;
wire net_3047;
wire net_16792;
wire net_8910;
wire net_9532;
wire net_6944;
wire net_6883;
wire net_2657;
wire net_15119;
wire net_12259;
wire net_11438;
wire net_14696;
wire net_8415;
wire net_7742;
wire net_2629;
wire net_2486;
wire net_15196;
wire net_7117;
wire net_16235;
wire net_1206;
wire net_8381;
wire net_3653;
wire x712;
wire net_13494;
wire net_1166;
wire net_17958;
wire net_18241;
wire net_10765;
wire net_801;
wire net_2620;
wire net_7450;
wire net_1718;
wire net_2581;
wire net_18318;
wire net_5093;
wire net_9417;
wire net_7372;
wire net_11921;
wire net_10391;
wire net_15612;
wire net_8482;
wire net_2129;
wire net_5968;
wire net_18131;
wire net_6234;
wire net_15112;
wire net_18896;
wire net_9833;
wire net_16156;
wire net_8856;
wire net_11382;
wire net_7115;
wire net_5906;
wire net_11391;
wire net_8462;
wire net_16797;
wire net_17412;
wire net_2325;
wire net_8807;
wire net_19011;
wire net_13715;
wire net_806;
wire net_11907;
wire net_9901;
wire net_16159;
wire net_18829;
wire net_18398;
wire net_16814;
wire net_8940;
wire net_4021;
wire net_17593;
wire net_10960;
wire net_946;
wire net_17156;
wire net_2194;
wire net_5010;
wire net_3559;
wire net_8370;
wire net_4682;
wire net_15261;
wire net_10114;
wire net_10402;
wire net_12499;
wire net_10732;
wire net_3564;
wire net_1448;
wire net_392;
wire net_5683;
wire net_7003;
wire net_2452;
wire net_11463;
wire net_10336;
wire net_3523;
wire net_4162;
wire net_17651;
wire net_5549;
wire net_3712;
wire net_6680;
wire x801;
wire net_16299;
wire net_17814;
wire net_1186;
wire net_4747;
wire net_14829;
wire net_7074;
wire net_17263;
wire net_10607;
wire net_10437;
wire net_2216;
wire net_10410;
wire net_16522;
wire net_7399;
wire net_3773;
wire net_1773;
wire net_9057;
wire net_8731;
wire net_18618;
wire net_17619;
wire net_5073;
wire net_4452;
wire net_2447;
wire net_7433;
wire net_14116;
wire net_5417;
wire net_15237;
wire net_8137;
wire net_14643;
wire net_17451;
wire net_182;
wire net_4359;
wire net_14506;
wire net_11260;
wire net_9547;
wire net_18051;
wire net_14872;
wire net_14237;
wire net_16581;
wire net_11442;
wire net_1435;
wire net_1370;
wire x13870;
wire net_9462;
wire net_3568;
wire net_4482;
wire net_6470;
wire net_19037;
wire net_8459;
wire net_1970;
wire net_1306;
wire net_1858;
wire net_14551;
wire x4059;
wire net_14846;
wire net_11332;
wire net_11196;
wire net_12242;
wire net_791;
wire net_14207;
wire net_9422;
wire net_1419;
wire net_3239;
wire net_8554;
wire net_2188;
wire net_17864;
wire net_12064;
wire net_13882;
wire net_17124;
wire net_17622;
wire net_14841;
wire net_7410;
wire net_12471;
wire net_7219;
wire net_13272;
wire net_6824;
wire net_14651;
wire net_361;
wire net_2890;
wire net_11547;
wire net_16991;
wire net_1905;
wire net_2540;
wire net_2230;
wire net_144;
wire net_227;
wire net_13758;
wire net_4183;
wire net_18368;
wire net_10237;
wire net_16788;
wire net_14664;
wire net_3592;
wire net_5961;
wire net_13728;
wire net_12543;
wire net_7156;
wire net_14413;
wire net_12636;
wire net_4969;
wire net_18926;
wire net_16817;
wire net_1415;
wire net_7052;
wire net_8859;
wire net_6379;
wire net_3317;
wire net_11746;
wire net_8140;
wire net_14934;
wire net_18531;
wire net_18162;
wire net_11638;
wire net_9161;
wire net_10120;
wire net_11910;
wire net_1230;
wire net_18126;
wire net_6047;
wire net_15418;
wire net_6862;
wire net_6064;
wire net_18204;
wire net_16850;
wire net_15455;
wire net_15317;
wire net_18577;
wire net_12046;
wire net_7585;
wire net_10597;
wire net_18138;
wire net_2039;
wire net_11579;
wire net_12067;
wire net_1456;
wire net_9198;
wire net_2227;
wire net_16822;
wire net_10280;
wire net_8876;
wire net_6968;
wire net_11041;
wire net_13509;
wire net_13844;
wire net_8752;
wire net_11209;
wire net_218;
wire net_12338;
wire net_16975;
wire net_7110;
wire net_9335;
wire net_5173;
wire net_1273;
wire net_3283;
wire net_18863;
wire net_9025;
wire net_4433;
wire net_17023;
wire net_13907;
wire net_11995;
wire net_2114;
wire net_2506;
wire net_5012;
wire net_9644;
wire net_16183;
wire net_7124;
wire net_18172;
wire net_11235;
wire net_11990;
wire net_16060;
wire net_14073;
wire net_285;
wire net_18078;
wire net_2499;
wire net_11567;
wire net_1297;
wire net_18822;
wire net_8901;
wire net_2177;
wire net_6581;
wire net_6916;
wire x4254;
wire net_16322;
wire net_18381;
wire net_17840;
wire net_5030;
wire net_1317;
wire net_215;
wire net_2394;
wire net_1382;
wire net_11593;
wire net_13408;
wire net_18171;
wire net_15513;
wire net_6442;
wire net_15487;
wire net_4508;
wire x13674;
wire net_17336;
wire net_8093;
wire net_3498;
wire net_12831;
wire net_13580;
wire net_9658;
wire net_5954;
wire net_14321;
wire net_6119;
wire net_14020;
wire net_9960;
wire net_16190;
wire net_14949;
wire net_10672;
wire net_16486;
wire net_10476;
wire net_16502;
wire net_2207;
wire net_263;
wire net_16027;
wire net_8509;
wire net_14139;
wire net_3483;
wire net_6838;
wire net_10548;
wire net_17936;
wire x170;
wire net_12528;
wire x725;
wire net_4189;
wire net_19034;
wire net_16826;
wire net_9256;
wire net_1090;
wire net_14850;
wire net_3685;
wire net_7030;
wire net_7012;
wire net_14107;
wire net_9007;
wire net_4285;
wire net_8643;
wire net_15862;
wire net_10726;
wire x52;
wire net_201;
wire net_5077;
wire net_17315;
wire net_9496;
wire x2068;
wire net_3280;
wire net_17426;
wire net_9666;
wire net_3085;
wire net_4043;
wire net_12631;
wire net_12207;
wire net_1852;
wire net_11236;
wire net_11912;
wire net_9515;
wire net_6129;
wire net_2780;
wire net_18631;
wire x608;
wire net_789;
wire net_15240;
wire net_10769;
wire net_3244;
wire net_12819;
wire net_9041;
wire net_15282;
wire net_18460;
wire net_12080;
wire net_3833;
wire net_9967;
wire net_8664;
wire net_7256;
wire net_14870;
wire net_8143;
wire net_5137;
wire net_17502;
wire net_11569;
wire net_1860;
wire net_18197;
wire net_14587;
wire net_8025;
wire net_1432;
wire net_1312;
wire net_9474;
wire net_5463;
wire net_16144;
wire net_8843;
wire net_8435;
wire net_4801;
wire net_16546;
wire net_5334;
wire net_16452;
wire net_5290;
wire net_14958;
wire net_17488;
wire net_3546;
wire net_8002;
wire net_1453;
wire net_14328;
wire net_13802;
wire net_13075;
wire net_9603;
wire net_3542;
wire net_634;
wire net_5374;
wire net_8516;
wire net_14177;
wire net_9630;
wire net_8055;
wire net_14066;
wire net_371;
wire net_15474;
wire net_13786;
wire net_7752;
wire net_2787;
wire net_2466;
wire net_4904;
wire net_8580;
wire net_4699;
wire net_7710;
wire net_7975;
wire net_8872;
wire net_18749;
wire net_7574;
wire net_13921;
wire net_18199;
wire net_5217;
wire net_17794;
wire net_679;
wire net_2680;
wire net_8116;
wire net_8924;
wire net_308;
wire net_12218;
wire net_6327;
wire net_890;
wire net_15693;
wire net_7228;
wire net_9019;
wire net_13401;
wire net_17269;
wire net_9162;
wire net_13646;
wire net_13595;
wire net_2471;
wire net_18643;
wire net_17524;
wire net_2404;
wire net_481;
wire net_16417;
wire net_5346;
wire net_18879;
wire net_16925;
wire net_6891;
wire net_11482;
wire net_1188;
wire net_13855;
wire net_1446;
wire net_541;
wire x9;
wire net_18309;
wire net_13380;
wire net_1251;
wire net_8157;
wire net_17725;
wire net_16301;
wire net_8830;
wire net_1697;
wire net_15748;
wire net_15741;
wire x13126;
wire net_4222;
wire net_12238;
wire net_1753;
wire net_4163;
wire net_14418;
wire net_5548;
wire net_14760;
wire net_14298;
wire net_4264;
wire net_9749;
wire net_18492;
wire net_17806;
wire net_15205;
wire net_9908;
wire net_11418;
wire net_7525;
wire net_17539;
wire net_3071;
wire net_8611;
wire net_14238;
wire net_10925;
wire net_9568;
wire net_7149;
wire net_9994;
wire net_7619;
wire net_16404;
wire net_2998;
wire x1532;
wire net_15549;
wire net_243;
wire net_8905;
wire net_6882;
wire net_2854;
wire net_10730;
wire net_17567;
wire net_8867;
wire net_4132;
wire net_8925;
wire net_4990;
wire net_7721;
wire net_9292;
wire net_16831;
wire net_11056;
wire net_13588;
wire net_8326;
wire net_1915;
wire net_17094;
wire net_15289;
wire net_13566;
wire net_10992;
wire net_8280;
wire net_18428;
wire net_4334;
wire net_16111;
wire net_14650;
wire net_17541;
wire net_15295;
wire net_18662;
wire net_12738;
wire net_18399;
wire net_13779;
wire net_12497;
wire net_18304;
wire net_18721;
wire net_14452;
wire net_18557;
wire net_17893;
wire net_13607;
wire net_15131;
wire net_17730;
wire net_9195;
wire net_17103;
wire net_12714;
wire net_7164;
wire net_12313;
wire net_14645;
wire net_9670;
wire net_14684;
wire net_7633;
wire net_13393;
wire net_18716;
wire net_17873;
wire net_8994;
wire net_3202;
wire net_13422;
wire net_4059;
wire net_6376;
wire net_6736;
wire net_7461;
wire net_15032;
wire net_15389;
wire net_10380;
wire net_5612;
wire net_2668;
wire net_13480;
wire net_2677;
wire net_15307;
wire net_14498;
wire net_15545;
wire net_10415;
wire net_11540;
wire net_11741;
wire net_3916;
wire net_6852;
wire net_8312;
wire net_13937;
wire net_18679;
wire net_14466;
wire net_12590;
wire net_18666;
wire net_5900;
wire net_6206;
wire net_3990;
wire net_10221;
wire net_3856;
wire net_9210;
wire net_17111;
wire net_17478;
wire net_5345;
wire net_8363;
wire net_4885;
wire net_17961;
wire net_14459;
wire net_3501;
wire net_16758;
wire net_7862;
wire net_12775;
wire net_6678;
wire net_15070;
wire net_7916;
wire net_13600;
wire net_8081;
wire x13567;
wire net_15524;
wire net_13982;
wire net_14013;
wire net_8835;
wire net_1272;
wire net_17743;
wire net_10273;
wire net_3505;
wire net_4001;
wire net_5059;
wire net_655;
wire net_3536;
wire net_6878;
wire net_16918;
wire net_8534;
wire net_10059;
wire net_17634;
wire net_18350;
wire net_16275;
wire net_12961;
wire net_9110;
wire net_14403;
wire net_423;
wire net_3036;
wire net_18446;
wire net_328;
wire net_10103;
wire net_10565;
wire net_7934;
wire net_7977;
wire net_9060;
wire net_3294;
wire net_3016;
wire net_4477;
wire net_12933;
wire net_9117;
wire net_11717;
wire net_3749;
wire net_2746;
wire net_12592;
wire net_9403;
wire net_5024;
wire net_15820;
wire net_18267;
wire net_14574;
wire net_11863;
wire net_2594;
wire net_15574;
wire net_17452;
wire net_17151;
wire net_5944;
wire net_15436;
wire net_811;
wire net_1684;
wire net_14549;
wire net_1462;
wire net_15019;
wire net_9150;
wire net_4993;
wire net_1926;
wire net_3115;
wire net_16621;
wire net_14158;
wire net_14809;
wire net_3518;
wire net_13069;
wire net_10261;
wire net_18335;
wire net_3680;
wire net_6926;
wire net_14319;
wire net_3984;
wire net_13317;
wire net_3615;
wire net_9559;
wire net_13172;
wire net_3055;
wire net_9844;
wire net_17813;
wire net_15782;
wire net_17230;
wire net_2845;
wire net_3095;
wire net_6510;
wire net_12585;
wire net_11358;
wire net_4586;
wire net_14986;
wire net_13141;
wire net_1763;
wire net_6168;
wire net_7291;
wire net_18338;
wire net_15476;
wire net_11067;
wire net_12999;
wire x1010;
wire net_3278;
wire net_12277;
wire net_4386;
wire net_8837;
wire net_1513;
wire net_15014;
wire net_16447;
wire net_10668;
wire net_12701;
wire net_4613;
wire net_7763;
wire net_11388;
wire net_10084;
wire net_3135;
wire net_5266;
wire net_5165;
wire net_8473;
wire net_18518;
wire net_8209;
wire net_1899;
wire net_15715;
wire net_8890;
wire net_4746;
wire net_16614;
wire net_12198;
wire net_1843;
wire net_6031;
wire net_17196;
wire net_12211;
wire net_7019;
wire net_534;
wire net_3793;
wire net_9261;
wire net_13523;
wire net_8659;
wire net_6823;
wire net_17316;
wire net_1551;
wire net_14951;
wire net_486;
wire net_18083;
wire net_14753;
wire net_12898;
wire net_406;
wire net_4190;
wire net_5391;
wire net_12448;
wire net_8967;
wire net_15186;
wire net_3640;
wire net_18455;
wire net_748;
wire net_10587;
wire net_6917;
wire net_13124;
wire net_10778;
wire net_3958;
wire net_12270;
wire net_5427;
wire net_16337;
wire net_15259;
wire net_11621;
wire net_11684;
wire net_14902;
wire net_514;
wire net_18766;
wire net_3645;
wire net_1604;
wire net_6499;
wire net_5755;
wire net_524;
wire net_13816;
wire net_17295;
wire net_4368;
wire net_7109;
wire net_13002;
wire net_18190;
wire net_3748;
wire net_15164;
wire net_10786;
wire net_9355;
wire net_14789;
wire net_12083;
wire net_5067;
wire net_10935;
wire net_1097;
wire net_11756;
wire net_12227;
wire net_14172;
wire net_762;
wire net_17176;
wire net_17373;
wire net_3589;
wire net_4943;
wire net_17766;
wire net_15827;
wire net_8400;
wire net_6173;
wire net_893;
wire net_3330;
wire net_11163;
wire net_255;
wire net_9641;
wire net_619;
wire net_13618;
wire net_9085;
wire net_17275;
wire net_3932;
wire net_7233;
wire net_11177;
wire net_7689;
wire net_14802;
wire net_7104;
wire net_14909;
wire net_3444;
wire net_4922;
wire net_3800;
wire net_3285;
wire net_17990;
wire net_7278;
wire net_4425;
wire net_18771;
wire net_4933;
wire net_5834;
wire net_17623;
wire net_4044;
wire net_14862;
wire net_11300;
wire net_13285;
wire net_11699;
wire net_5875;
wire net_4630;
wire net_16091;
wire net_15636;
wire net_976;
wire net_6287;
wire net_2709;
wire net_5309;
wire net_10321;
wire net_11630;
wire net_611;
wire x4011;
wire net_7879;
wire net_17849;
wire net_3514;
wire net_5441;
wire net_17560;
wire net_6077;
wire net_10849;
wire net_4907;
wire net_6567;
wire net_4107;
wire net_18285;
wire net_2160;
wire net_3692;
wire net_3477;
wire net_391;
wire net_6361;
wire net_9268;
wire net_9723;
wire net_5040;
wire net_18108;
wire net_5820;
wire net_6692;
wire net_4172;
wire net_16735;
wire net_13892;
wire net_8123;
wire net_12417;
wire net_1141;
wire net_6253;
wire net_10621;
wire net_16372;
wire net_3243;
wire net_4867;
wire net_7871;
wire net_2104;
wire net_5564;
wire net_17040;
wire net_6190;
wire net_2766;
wire net_3771;
wire net_12469;
wire net_2417;
wire net_16004;
wire net_14406;
wire net_741;
wire x225;
wire net_5509;
wire net_17862;
wire net_15092;
wire net_7853;
wire net_6472;
wire net_13765;
wire net_3789;
wire net_15664;
wire net_13288;
wire net_18783;
wire net_9598;
wire net_11947;
wire net_12977;
wire net_2850;
wire net_770;
wire net_13905;
wire net_12901;
wire net_1005;
wire net_15711;
wire net_11792;
wire net_11198;
wire net_1059;
wire net_3891;
wire net_4918;
wire net_16650;
wire net_18903;
wire net_17240;
wire net_1796;
wire net_10328;
wire x2594;
wire net_5187;
wire net_7501;
wire net_11368;
wire net_11291;
wire net_1507;
wire net_2310;
wire net_18354;
wire net_7466;
wire net_474;
wire net_16901;
wire net_16358;
wire net_12518;
wire net_11421;
wire net_11934;
wire net_18076;
wire net_11940;
wire net_7947;
wire net_16310;
wire net_11855;
wire net_12244;
wire net_944;
wire net_16019;
wire net_10008;
wire net_17385;
wire net_18236;
wire net_13477;
wire net_12538;
wire net_11002;
wire net_7199;
wire net_12580;
wire net_17003;
wire net_15709;
wire net_13669;
wire net_12028;
wire net_287;
wire net_17492;
wire net_189;
wire net_10414;
wire net_9893;
wire net_9860;
wire net_15988;
wire net_3755;
wire net_6036;
wire net_433;
wire net_11709;
wire net_8296;
wire net_4443;
wire net_224;
wire net_15886;
wire net_1898;
wire net_9073;
wire net_608;
wire net_1212;
wire net_3604;
wire net_4383;
wire net_5331;
wire net_13194;
wire net_3706;
wire net_16387;
wire net_7062;
wire net_12879;
wire net_11997;
wire net_8299;
wire net_12832;
wire net_18066;
wire net_18443;
wire net_6416;
wire net_16696;
wire net_15923;
wire net_13227;
wire net_17573;
wire net_873;
wire net_1811;
wire net_13884;
wire net_12374;
wire net_11080;
wire net_2588;
wire net_7802;
wire net_18921;
wire net_9771;
wire net_704;
wire net_12906;
wire net_3997;
wire net_1356;
wire net_14542;
wire net_8913;
wire net_4393;
wire net_6541;
wire net_3816;
wire net_6101;
wire net_13457;
wire net_5539;
wire net_9056;
wire net_1711;
wire net_14527;
wire net_2084;
wire net_8186;
wire net_11590;
wire net_9530;
wire net_5085;
wire net_7031;
wire net_7349;
wire net_12653;
wire net_8680;
wire net_16506;
wire net_4836;
wire net_9602;
wire net_17366;
wire net_15265;
wire net_11663;
wire net_7270;
wire net_9283;
wire net_12892;
wire net_2526;
wire net_18758;
wire net_16237;
wire net_9414;
wire net_18838;
wire net_7338;
wire net_1644;
wire net_12126;
wire net_2800;
wire net_14225;
wire net_7940;
wire net_17354;
wire net_17695;
wire net_8255;
wire net_1190;
wire net_3225;
wire net_4093;
wire net_6449;
wire net_15535;
wire net_4799;
wire net_16269;
wire net_13812;
wire net_8721;
wire net_12021;
wire net_9829;
wire net_6066;
wire net_17361;
wire net_15140;
wire net_2191;
wire net_14698;
wire net_13318;
wire net_13304;
wire net_10690;
wire x1885;
wire net_17672;
wire net_15077;
wire net_13168;
wire net_12617;
wire net_15639;
wire net_12416;
wire net_12352;
wire net_14249;
wire net_1577;
wire net_17714;
wire net_1054;
wire net_4595;
wire net_17595;
wire net_2727;
wire net_18225;
wire net_16185;
wire net_5605;
wire net_2257;
wire net_10640;
wire net_14741;
wire net_3418;
wire net_18751;
wire net_5491;
wire net_13217;
wire net_12044;
wire net_2968;
wire net_7314;
wire net_10649;
wire net_5989;
wire net_16105;
wire net_12339;
wire net_2643;
wire net_5845;
wire net_9591;
wire net_3722;
wire net_18034;
wire net_11117;
wire net_17739;
wire net_18331;
wire net_1517;
wire net_16416;
wire net_11218;
wire net_5980;
wire net_6705;
wire net_9192;
wire net_15217;
wire net_1690;
wire net_16606;
wire net_11924;
wire net_2093;
wire net_2997;
wire net_14831;
wire net_15027;
wire net_14186;
wire net_9076;
wire net_7239;
wire net_18776;
wire net_11787;
wire net_17138;
wire net_15099;
wire net_18419;
wire net_9549;
wire net_4357;
wire net_16878;
wire net_16714;
wire net_2536;
wire net_5890;
wire net_7968;
wire x13488;
wire x1281;
wire net_2949;
wire net_3429;
wire net_10954;
wire net_9032;
wire net_1708;
wire net_12398;
wire net_5519;
wire net_17215;
wire net_15966;
wire net_13112;
wire net_12575;
wire net_13050;
wire net_722;
wire net_5420;
wire net_17065;
wire net_12094;
wire net_18044;
wire net_14612;
wire net_13099;
wire net_5798;
wire net_11351;
wire net_14313;
wire net_5223;
wire net_8216;
wire net_435;
wire net_12077;
wire net_1830;
wire net_5156;
wire net_6481;
wire net_1649;
wire net_6603;
wire net_1837;
wire net_6973;
wire net_2427;
wire net_8075;
wire net_1071;
wire net_3378;
wire net_18607;
wire net_5004;
wire net_5817;
wire net_9776;
wire net_18499;
wire net_1701;
wire net_5675;
wire net_11156;
wire net_14007;
wire net_8678;
wire net_12175;
wire net_1633;
wire net_11132;
wire net_12150;
wire net_5251;
wire net_8694;
wire net_15759;
wire net_319;
wire net_18435;
wire net_2670;
wire net_1743;
wire net_2597;
wire net_5913;
wire net_7640;
wire net_11887;
wire net_4139;
wire net_2923;
wire net_7545;
wire net_512;
wire net_16646;
wire net_17878;
wire net_3102;
wire net_18027;
wire net_7510;
wire net_16221;
wire net_13513;
wire net_5780;
wire net_5721;
wire net_7904;
wire net_13119;
wire net_16368;
wire net_16243;
wire net_16999;
wire net_3371;
wire net_17898;
wire net_5317;
wire net_13953;
wire net_15874;
wire x1383;
wire net_6800;
wire net_9375;
wire net_12673;
wire net_17143;
wire net_15212;
wire net_1875;
wire net_5862;
wire net_3420;
wire net_3887;
wire net_18009;
wire net_16964;
wire net_7050;
wire x13853;
wire net_7484;
wire net_13373;
wire net_15045;
wire net_12189;
wire net_8736;
wire net_16585;
wire net_12953;
wire net_5178;
wire net_17035;
wire net_7678;
wire net_17463;
wire net_2835;
wire net_4543;
wire net_4871;
wire net_6599;
wire net_1240;
wire net_9213;
wire net_3000;
wire net_16761;
wire net_12200;
wire net_15002;
wire net_15768;
wire net_12674;
wire net_17533;
wire net_13048;
wire net_858;
wire net_9338;
wire net_15583;
wire net_8986;
wire net_4766;
wire net_6004;
wire net_16167;
wire net_8504;
wire net_13549;
wire net_9867;
wire net_7995;
wire net_3735;
wire net_10870;
wire net_11422;
wire net_1427;
wire net_5123;
wire net_17980;
wire net_3921;
wire net_7075;
wire net_5899;
wire net_4098;
wire net_5478;
wire net_7251;
wire net_16494;
wire net_12106;
wire net_9827;
wire net_11029;
wire net_18676;
wire net_17702;
wire net_14762;
wire net_10308;
wire net_6020;
wire net_7172;
wire net_1677;
wire net_13260;
wire net_7089;
wire net_2811;
wire net_6788;
wire net_2612;
wire net_8791;
wire net_5230;
wire net_2042;
wire net_7189;
wire net_13626;
wire net_17218;
wire net_11649;
wire net_18270;
wire net_6649;
wire net_10949;
wire net_3488;
wire net_3023;
wire net_17010;
wire net_5584;
wire net_1202;
wire net_14373;
wire net_10890;
wire net_925;
wire net_4932;
wire net_6776;
wire net_7452;
wire net_12827;
wire net_5384;
wire net_17250;
wire net_15680;
wire net_11317;
wire net_10974;
wire net_12074;
wire net_4661;
wire net_2695;
wire net_10196;
wire net_11054;
wire net_14337;
wire net_13336;
wire net_12851;
wire net_12611;
wire net_7404;
wire net_8564;
wire net_7783;
wire net_14477;
wire net_18107;
wire net_6284;
wire net_9436;
wire net_7132;
wire net_2313;
wire net_11655;
wire net_9044;
wire net_6172;
wire net_7595;
wire net_230;
wire net_18472;
wire net_4214;
wire net_18861;
wire net_6985;
wire net_3349;
wire net_4782;
wire net_1222;
wire net_3404;
wire net_14080;
wire net_14291;
wire net_17734;
wire net_3810;
wire net_14560;
wire net_9172;
wire net_12018;
wire net_15689;
wire net_4739;
wire net_4156;
wire net_8823;
wire net_12685;
wire net_13693;
wire net_12459;
wire net_3440;
wire net_6904;
wire net_3358;
wire net_1776;
wire net_3368;
wire net_5747;
wire net_15897;
wire net_4014;
wire net_14723;
wire net_15626;
wire net_18116;
wire net_7204;
wire net_17017;
wire net_2132;
wire net_2292;
wire net_9313;
wire net_12367;
wire net_1880;
wire net_17856;
wire net_3862;
wire net_184;
wire net_5103;
wire net_17901;
wire net_5855;
wire net_10757;
wire net_14087;
wire net_11247;
wire net_10427;
wire net_15359;
wire net_7203;
wire net_18214;
wire net_18967;
wire net_17089;
wire net_1867;
wire net_18626;
wire net_9498;
wire net_8205;
wire net_1949;
wire net_2650;
wire net_13568;
wire net_10455;
wire net_1804;
wire net_17554;
wire net_2331;
wire net_14520;
wire net_6667;
wire net_16741;
wire net_16042;
wire net_4291;
wire net_12389;
wire net_8637;
wire net_14483;
wire net_1135;
wire net_1365;
wire net_16768;
wire net_11674;
wire net_1346;
wire net_5047;
wire net_18957;
wire net_17199;
wire net_11478;
wire net_15946;
wire net_13865;
wire net_13835;
wire net_9220;
wire net_9277;
wire net_1801;
wire net_18819;
wire net_15650;
wire net_14364;
wire net_4350;
wire net_6029;
wire net_8955;
wire net_15724;
wire net_669;
wire net_937;
wire net_11252;
wire net_10179;
wire net_8452;
wire net_9575;
wire net_8030;
wire net_479;
wire net_8740;
wire net_12769;
wire net_6086;
wire net_2030;
wire net_1587;
wire net_17077;
wire net_13232;
wire net_11025;
wire net_796;
wire net_18610;
wire net_648;
wire net_11901;
wire net_16109;
wire net_6884;
wire net_12040;
wire net_8150;
wire net_16888;
wire net_14300;
wire net_14443;
wire net_7054;
wire net_11950;
wire net_7625;
wire net_3658;
wire net_12560;
wire x4701;
wire net_14146;
wire net_6964;
wire net_9148;
wire net_15871;
wire net_15414;
wire net_18550;
wire net_17953;
wire net_8237;
wire net_17951;
wire net_17123;
wire net_8556;
wire net_7649;
wire net_16793;
wire net_15804;
wire net_12179;
wire net_10739;
wire net_10232;
wire net_15840;
wire net_8725;
wire net_4492;
wire net_6700;
wire net_14655;
wire net_1961;
wire net_10831;
wire net_1260;
wire net_10124;
wire net_9832;
wire net_15375;
wire net_239;
wire net_18824;
wire net_13396;
wire net_310;
wire net_18899;
wire net_14599;
wire net_10367;
wire net_2437;
wire net_10792;
wire net_14772;
wire net_8982;
wire net_9917;
wire net_13498;
wire net_5886;
wire net_14960;
wire net_17755;
wire net_13711;
wire net_682;
wire net_17580;
wire net_1963;
wire net_7122;
wire net_17114;
wire net_13558;
wire net_16033;
wire net_12049;
wire net_17976;
wire net_8989;
wire net_3560;
wire net_5804;
wire net_17908;
wire net_1007;
wire net_15497;
wire net_7000;
wire net_14837;
wire net_4772;
wire net_7007;
wire net_11415;
wire net_1292;
wire net_7197;
wire net_10703;
wire net_7861;
wire net_10771;
wire net_12262;
wire net_11039;
wire net_2796;
wire net_18202;
wire net_11400;
wire net_16526;
wire net_15845;
wire net_19044;
wire net_5016;
wire net_4024;
wire net_6699;
wire net_9544;
wire net_12443;
wire net_6280;
wire net_17086;
wire net_8043;
wire net_1937;
wire net_15114;
wire net_7215;
wire net_18308;
wire net_1956;
wire net_11339;
wire net_13433;
wire net_1614;
wire net_13491;
wire net_12911;
wire net_11958;
wire net_16597;
wire net_7119;
wire x13527;
wire net_10255;
wire net_3209;
wire net_12791;
wire net_4891;
wire net_8688;
wire net_10874;
wire net_8412;
wire net_7716;
wire net_294;
wire net_17606;
wire net_15305;
wire x563;
wire net_9837;
wire net_10797;
wire net_2429;
wire net_9217;
wire net_1265;
wire net_10822;
wire net_6224;
wire net_14694;
wire net_8697;
wire net_11203;
wire net_12984;
wire net_8039;
wire net_1619;
wire net_5468;
wire net_12727;
wire net_18742;
wire net_2124;
wire net_5934;
wire net_15247;
wire net_1161;
wire net_7070;
wire net_4671;
wire net_17587;
wire net_13606;
wire net_12695;
wire net_7663;
wire net_11385;
wire net_10721;
wire net_8500;
wire net_1395;
wire net_8877;
wire net_9360;
wire net_15005;
wire net_11875;
wire net_17128;
wire net_14678;
wire net_5353;
wire net_16195;
wire net_8756;
wire net_5270;
wire net_9921;
wire net_12456;
wire net_18218;
wire net_2445;
wire net_3396;
wire net_6640;
wire net_5324;
wire net_15452;
wire net_10592;
wire net_16836;
wire net_4511;
wire net_7395;
wire net_13419;
wire net_2894;
wire net_15643;
wire net_13714;
wire net_6999;
wire net_1988;
wire net_7388;
wire net_3718;
wire net_4419;
wire net_15619;
wire net_5284;
wire net_16488;
wire net_11125;
wire net_3525;
wire net_10696;
wire net_6850;
wire net_13508;
wire net_1608;
wire net_506;
wire net_3769;
wire net_12802;
wire net_8019;
wire net_9330;
wire net_12836;
wire net_3775;
wire net_8278;
wire net_5432;
wire net_6586;
wire net_5096;
wire net_16020;
wire x13011;
wire net_7589;
wire net_12055;
wire net_6909;
wire net_290;
wire net_6476;
wire net_13676;
wire net_6315;
wire net_10913;
wire net_3313;
wire net_9987;
wire net_8803;
wire net_5769;
wire net_3591;
wire net_5729;
wire net_16812;
wire net_16207;
wire net_13341;
wire net_15025;
wire net_16464;
wire net_11926;
wire net_12430;
wire net_4436;
wire net_15775;
wire net_2329;
wire net_16801;
wire net_2150;
wire net_7129;
wire net_2065;
wire net_10003;
wire net_13244;
wire net_10030;
wire net_17467;
wire net_8373;
wire net_2927;
wire net_7397;
wire net_16634;
wire net_11831;
wire net_11838;
wire net_194;
wire net_4856;
wire net_13941;
wire net_11264;
wire net_9448;
wire net_1128;
wire net_2713;
wire net_13161;
wire net_11582;
wire net_15354;
wire net_12539;
wire net_11320;
wire net_1119;
wire net_9637;
wire net_4312;
wire net_5299;
wire net_8852;
wire net_3345;
wire net_18319;
wire net_10125;
wire net_18582;
wire net_7855;
wire net_11642;
wire net_11006;
wire net_7127;
wire net_7448;
wire net_11900;
wire net_18042;
wire net_10742;
wire net_3328;
wire net_14812;
wire net_10174;
wire net_16328;
wire net_2107;
wire net_180;
wire net_13462;
wire net_17107;
wire net_6859;
wire net_5657;
wire net_4367;
wire net_3290;
wire net_3731;
wire net_1475;
wire net_10241;
wire net_18207;
wire net_14112;
wire net_16459;
wire net_16738;
wire net_10601;
wire net_5446;
wire net_12719;
wire net_2173;
wire net_18597;
wire net_9053;
wire net_6865;
wire net_7539;
wire net_14785;
wire net_6263;
wire net_5590;
wire net_11673;
wire net_14334;
wire net_5476;
wire net_3744;
wire net_11851;
wire net_4635;
wire net_14912;
wire net_12193;
wire net_18946;
wire net_6570;
wire net_8309;
wire net_15360;
wire net_6939;
wire net_12968;
wire net_4485;
wire net_1558;
wire net_8603;
wire net_4641;
wire net_17405;
wire net_10958;
wire net_10806;
wire net_14138;
wire net_455;
wire net_11515;
wire net_16072;
wire net_10294;
wire net_7498;
wire net_3339;
wire net_6303;
wire net_9428;
wire net_7352;
wire net_1832;
wire net_12474;
wire net_12622;
wire net_1026;
wire net_16095;
wire net_2215;
wire net_15376;
wire net_6453;
wire net_2573;
wire x2805;
wire net_9369;
wire net_10312;
wire x13474;
wire net_7378;
wire net_19004;
wire net_3993;
wire net_13673;
wire net_1401;
wire net_3909;
wire net_11858;
wire net_17800;
wire net_7889;
wire net_14394;
wire net_7248;
wire x3604;
wire net_13311;
wire net_17557;
wire net_443;
wire net_6367;
wire net_6495;
wire net_18907;
wire net_8486;
wire net_17661;
wire net_18389;
wire net_12364;
wire net_7956;
wire net_14034;
wire net_11346;
wire net_1990;
wire net_7456;
wire net_18155;
wire net_10442;
wire net_17350;
wire net_16391;
wire net_9951;
wire net_18843;
wire net_7880;
wire net_11988;
wire net_11601;
wire net_622;
wire net_17028;
wire net_14854;
wire net_11993;
wire net_11277;
wire net_5909;
wire net_11225;
wire net_1338;
wire net_7842;
wire net_2053;
wire net_6623;
wire net_2180;
wire net_4242;
wire net_2119;
wire net_3220;
wire net_4720;
wire net_18152;
wire net_13108;
wire net_8627;
wire net_7474;
wire net_5920;
wire net_6124;
wire net_8384;
wire net_6992;
wire net_13519;
wire net_2007;
wire net_5143;
wire net_5763;
wire net_7703;
wire net_16211;
wire net_713;
wire net_10653;
wire net_5711;
wire net_17329;
wire net_16898;
wire net_13338;
wire net_8700;
wire net_11104;
wire net_729;
wire net_9222;
wire net_4197;
wire net_17292;
wire net_14893;
wire net_13156;
wire net_7093;
wire net_7324;
wire net_13948;
wire net_9169;
wire net_8447;
wire net_5366;
wire net_14596;
wire net_8711;
wire net_13571;
wire net_341;
wire net_13611;
wire net_14733;
wire net_12992;
wire net_970;
wire net_13362;
wire net_13389;
wire net_8653;
wire net_15539;
wire net_15984;
wire net_13917;
wire net_13184;
wire net_3044;
wire net_5929;
wire net_17257;
wire net_17457;
wire net_11145;
wire net_14745;
wire net_13726;
wire net_14071;
wire net_14233;
wire net_12038;
wire net_10100;
wire net_2163;
wire net_3417;
wire x4234;
wire net_3307;
wire net_13301;
wire net_12534;
wire net_553;
wire net_4212;
wire net_6133;
wire net_7797;
wire net_8300;
wire net_6239;
wire net_15991;
wire net_4701;
wire net_18262;
wire net_10889;
wire net_15906;
wire net_462;
wire net_418;
wire net_15415;
wire net_15105;
wire net_161;
wire net_7988;
wire net_17615;
wire net_8660;
wire net_1486;
wire net_2606;
wire net_18687;
wire net_1839;
wire net_2320;
wire net_1665;
wire net_11076;
wire net_14515;
wire net_13744;
wire net_8525;
wire net_8349;
wire net_18900;
wire net_16179;
wire net_3550;
wire net_16663;
wire net_12377;
wire net_11172;
wire net_16056;
wire net_6893;
wire net_9466;
wire net_2224;
wire net_7066;
wire net_10037;
wire net_15404;
wire net_5733;
wire net_15847;
wire net_2458;
wire net_9324;
wire net_17164;
wire net_3435;
wire net_2635;
wire net_16789;
wire net_3374;
wire net_5207;
wire net_15490;
wire net_13540;
wire net_5572;
wire net_15068;
wire net_8283;
wire net_1037;
wire net_2019;
wire net_18379;
wire net_4676;
wire net_8395;
wire net_6675;
wire net_13033;
wire net_7549;
wire net_6793;
wire net_15793;
wire x735;
wire net_17668;
wire net_6242;
wire net_14433;
wire net_15012;
wire net_1623;
wire net_2982;
wire net_6948;
wire net_4410;
wire net_7230;
wire net_16849;
wire net_5785;
wire net_14047;
wire net_18245;
wire net_17514;
wire net_18537;
wire net_14251;
wire net_13657;
wire net_8650;
wire net_7190;
wire net_10907;
wire net_16000;
wire net_18299;
wire net_8596;
wire net_10984;
wire net_12147;
wire net_12166;
wire net_6651;
wire net_16009;
wire net_5485;
wire net_7243;
wire net_18974;
wire net_12004;
wire net_3554;
wire net_12323;
wire net_1920;
wire net_4101;
wire net_17628;
wire net_2010;
wire net_18913;
wire net_11665;
wire net_8782;
wire net_6941;
wire net_8321;
wire net_9139;
wire net_16853;
wire net_18507;
wire net_4672;
wire net_8862;
wire net_6743;
wire net_1723;
wire net_8465;
wire net_2900;
wire net_14790;
wire net_17648;
wire net_11015;
wire net_5152;
wire net_5718;
wire net_8190;
wire net_17396;
wire net_4376;
wire net_17288;
wire net_14397;
wire net_18881;
wire net_16868;
wire net_2306;
wire net_12382;
wire net_2873;
wire net_3272;
wire net_14618;
wire net_2254;
wire net_2861;
wire net_18235;
wire net_11844;
wire net_14343;
wire net_9570;
wire net_4574;
wire net_18701;
wire net_1209;
wire net_15936;
wire net_13076;
wire net_4038;
wire net_847;
wire net_10157;
wire net_4787;
wire net_11740;
wire net_283;
wire net_12864;
wire net_13505;
wire net_5117;
wire net_18875;
wire net_4690;
wire net_12796;
wire net_5020;
wire net_14126;
wire net_7316;
wire net_5445;
wire net_18725;
wire net_7428;
wire net_10023;
wire net_10990;
wire net_7958;
wire net_16559;
wire net_344;
wire net_14102;
wire net_4757;
wire net_18735;
wire net_15956;
wire net_2269;
wire net_884;
wire net_14184;
wire net_712;
wire net_1422;
wire net_2281;
wire net_12940;
wire net_17655;
wire net_4497;
wire net_11527;
wire net_18960;
wire net_6670;
wire net_15061;
wire net_1106;
wire net_15817;
wire net_13629;
wire net_8483;
wire net_2972;
wire net_5611;
wire net_11311;
wire net_10836;
wire net_15252;
wire net_2241;
wire net_13006;
wire net_17430;
wire net_9522;
wire net_8615;
wire net_1547;
wire net_15596;
wire net_13053;
wire net_8768;
wire net_5122;
wire net_12495;
wire net_11146;
wire net_5423;
wire net_13972;
wire x1690;
wire net_7971;
wire net_6507;
wire net_9912;
wire net_10395;
wire net_7344;
wire net_16956;
wire net_5055;
wire net_14886;
wire net_7303;
wire net_17392;
wire net_4794;
wire net_2625;
wire net_4149;
wire net_5687;
wire net_6849;
wire net_10292;
wire x641;
wire net_1595;
wire net_5849;
wire net_15656;
wire net_12919;
wire x2261;
wire net_3432;
wire net_2974;
wire net_6519;
wire net_14517;
wire net_3895;
wire net_8339;
wire net_13660;
wire net_11736;
wire net_2734;
wire net_12888;
wire net_18603;
wire net_15508;
wire net_13133;
wire net_10637;
wire net_12569;
wire net_6761;
wire net_14857;
wire net_3146;
wire net_6294;
wire net_7827;
wire net_18118;
wire net_6390;
wire net_9347;
wire net_10496;
wire net_5237;
wire net_16601;
wire net_14825;
wire net_17643;
wire net_11553;
wire net_3022;
wire net_8226;
wire net_10989;
wire net_16808;
wire net_7495;
wire net_9616;
wire net_5741;
wire net_6391;
wire net_8476;
wire net_6308;
wire net_18513;
wire net_16170;
wire x4561;
wire net_17344;
wire net_5700;
wire net_7441;
wire net_9671;
wire net_15405;
wire net_9159;
wire net_11899;
wire net_14260;
wire net_18684;
wire net_18473;
wire net_4706;
wire net_594;
wire net_5532;
wire net_17203;
wire net_11336;
wire net_9818;
wire net_17225;
wire net_14310;
wire net_11892;
wire net_8512;
wire net_11690;
wire net_6188;
wire net_4402;
wire net_6328;
wire net_2074;
wire net_16254;
wire net_8428;
wire net_5256;
wire net_16842;
wire net_5274;
wire net_10183;
wire net_2577;
wire net_11091;
wire net_8286;
wire net_2954;
wire net_15890;
wire net_3274;
wire net_17762;
wire net_16143;
wire net_2953;
wire net_15731;
wire net_6380;
wire net_467;
wire net_2910;
wire net_8728;
wire net_4851;
wire net_2081;
wire net_9245;
wire net_10522;
wire net_5195;
wire net_11426;
wire net_18132;
wire net_14555;
wire net_3165;
wire net_12644;
wire net_18858;
wire net_4965;
wire net_12295;
wire net_8648;
wire net_2302;
wire net_12523;
wire net_18280;
wire net_14601;
wire net_8545;
wire net_13649;
wire net_5502;
wire net_6805;
wire net_6387;
wire net_6403;
wire net_7734;
wire net_18344;
wire net_13873;
wire net_12409;
wire net_15916;
wire net_15294;
wire net_2368;
wire net_18482;
wire net_19001;
wire net_12908;
wire net_3966;
wire net_6330;
wire net_607;
wire net_12392;
wire net_8106;
wire net_9739;
wire net_4142;
wire net_1045;
wire net_3497;
wire net_3905;
wire net_13087;
wire net_15392;
wire net_13249;
wire net_4939;
wire x13501;
wire net_17246;
wire net_3601;
wire net_9933;
wire net_16133;
wire net_4538;
wire net_19041;
wire net_14648;
wire net_13044;
wire net_12052;
wire net_18073;
wire net_15550;
wire net_11167;
wire net_16685;
wire net_12662;
wire net_4527;
wire net_6419;
wire net_18187;
wire net_8548;
wire net_4144;
wire net_4716;
wire net_7586;
wire net_2079;
wire net_1731;
wire net_2052;
wire net_16038;
wire net_9089;
wire net_16541;
wire net_9648;
wire net_9463;
wire net_6912;
wire net_12813;
wire net_17419;
wire net_13276;
wire net_17202;
wire net_5952;
wire net_11769;
wire net_15422;
wire net_3636;
wire net_7184;
wire net_14095;
wire net_4727;
wire net_17769;
wire net_5032;
wire net_11046;
wire net_1536;
wire net_5852;
wire net_6232;
wire net_12504;
wire net_3478;
wire net_1498;
wire net_8117;
wire net_18089;
wire net_10815;
wire net_5561;
wire net_5626;
wire net_949;
wire net_14000;
wire net_12401;
wire net_10936;
wire net_7813;
wire net_4111;
wire net_9392;
wire net_14267;
wire net_10616;
wire net_12947;
wire net_12287;
wire net_18359;
wire net_18141;
wire net_12722;
wire net_14283;
wire net_8262;
wire net_9028;
wire net_2296;
wire net_9438;
wire net_13994;
wire net_3385;
wire net_17798;
wire net_357;
wire net_6954;
wire net_9179;
wire net_12934;
wire net_7849;
wire net_3451;
wire net_18769;
wire net_7085;
wire net_8790;
wire net_2694;
wire net_17184;
wire net_12280;
wire net_5607;
wire net_2096;
wire net_3118;
wire net_5555;
wire net_18560;
wire net_18521;
wire net_15330;
wire net_11501;
wire net_1829;
wire net_16434;
wire net_14240;
wire net_13904;
wire x13403;
wire net_9780;
wire net_662;
wire net_862;
wire net_16121;
wire net_2307;
wire net_7168;
wire net_14822;
wire net_8127;
wire net_4174;
wire net_5396;
wire net_738;
wire net_4080;
wire net_4325;
wire net_1150;
wire net_504;
wire net_18831;
wire net_10333;
wire net_9789;
wire x3712;
wire net_6634;
wire net_11537;
wire net_7698;
wire net_17839;
wire net_16593;
wire net_18348;
wire net_3120;
wire net_14324;
wire net_18274;
wire net_4504;
wire net_1561;
wire net_12161;
wire net_3269;
wire net_11455;
wire net_17332;
wire net_10472;
wire net_4421;
wire net_18360;
wire net_6666;
wire net_17048;
wire net_17775;
wire net_13329;
wire net_9855;
wire net_1940;
wire net_13323;
wire net_11449;
wire net_10452;
wire net_8635;
wire net_11516;
wire x14005;
wire net_16670;
wire net_12781;
wire net_14621;
wire net_11528;
wire net_991;
wire net_3912;
wire net_6528;
wire net_13204;
wire net_18253;
wire net_6753;
wire net_3088;
wire net_11107;
wire net_4607;
wire net_12484;
wire net_2979;
wire net_17925;
wire net_16712;
wire net_10714;
wire net_2772;
wire x4831;
wire net_9564;
wire net_8491;
wire net_5775;
wire net_4180;
wire net_15562;
wire net_13839;
wire net_12116;
wire net_12180;
wire net_2347;
wire net_11710;
wire net_14777;
wire net_2684;
wire net_3806;
wire net_10795;
wire net_10352;
wire net_521;
wire net_3972;
wire net_14275;
wire net_9003;
wire net_14738;
wire net_2754;
wire net_267;
wire net_1585;
wire net_13748;
wire net_11613;
wire net_9143;
wire net_18541;
wire net_11099;
wire net_15761;
wire net_6898;
wire net_7421;
wire net_16618;
wire net_3663;
wire net_10885;
wire net_3260;
wire net_5110;
wire net_13017;
wire net_9186;
wire net_6465;
wire net_6486;
wire net_6048;
wire net_13177;
wire net_18652;
wire net_2716;
wire net_11815;
wire net_6551;
wire net_4750;
wire net_15868;
wire net_13346;
wire net_4558;
wire net_12858;
wire x468;
wire net_8394;
wire net_15521;
wire net_2828;
wire net_12749;
wire net_824;
wire net_3458;
wire net_1822;
wire net_18801;
wire net_9755;
wire net_13038;
wire net_1972;
wire net_15559;
wire x4635;
wire net_17945;
wire net_12267;
wire net_3126;
wire net_993;
wire net_10555;
wire net_5974;
wire net_9456;
wire net_1100;
wire net_7035;
wire net_15121;
wire net_14995;
wire net_2817;
wire net_18039;
wire net_6686;
wire net_10046;
wire net_17931;
wire net_15128;
wire x3925;
wire net_5996;
wire net_6730;
wire net_13823;
wire net_1326;
wire net_7488;
wire net_546;
wire net_4648;
wire net_14638;
wire net_4546;
wire net_10065;
wire net_13735;
wire net_13320;
wire net_8062;
wire net_17987;
wire net_12424;
wire net_3701;
wire net_18712;
wire net_17147;
wire net_14296;
wire net_4736;
wire net_7592;
wire net_5592;
wire net_5642;
wire net_8012;
wire net_7906;
wire net_4974;
wire net_3883;
wire net_1542;
wire net_17546;
wire net_1172;
wire x4964;
wire net_9124;
wire net_13703;
wire net_8431;
wire net_4230;
wire net_14626;
wire net_16747;
wire net_16228;
wire net_9503;
wire net_4860;
wire net_2237;
wire net_2566;
wire net_8352;
wire net_3953;
wire net_917;
wire net_3730;
wire net_2874;
wire net_10965;
wire net_8942;
wire net_14535;
wire net_9685;
wire net_2993;
wire net_18146;
wire net_10921;
wire net_3067;
wire net_13950;
wire net_10075;
wire net_4288;
wire x13969;
wire net_323;
wire net_5402;
wire net_963;
wire net_10301;
wire net_16534;
wire net_9482;
wire net_7368;
wire net_4689;
wire net_10216;
wire net_153;
wire net_2389;
wire net_12328;
wire net_6276;
wire net_7556;
wire net_375;
wire net_562;
wire net_16692;
wire net_364;
wire net_8675;
wire net_14380;
wire net_12770;
wire net_17802;
wire net_11723;
wire net_3172;
wire net_10485;
wire net_13772;
wire net_11706;
wire net_4239;
wire net_14011;
wire net_5516;
wire net_7177;
wire net_6313;
wire net_16535;
wire net_6341;
wire net_8161;
wire net_6840;
wire net_18111;
wire net_12810;
wire net_18567;
wire net_3171;
wire net_7514;
wire net_14217;
wire net_12742;
wire net_17511;
wire net_14472;
wire net_10091;
wire net_8173;
wire net_1247;
wire net_3673;
wire net_18793;
wire net_11149;
wire net_2388;
wire net_15383;
wire net_14006;
wire net_16396;
wire net_1215;
wire net_5169;
wire net_5248;
wire net_15578;
wire x3122;
wire net_284;
wire net_6655;
wire net_12743;
wire net_439;
wire net_18322;
wire net_259;
wire net_3582;
wire net_3351;
wire net_4094;
wire net_18977;
wire net_18505;
wire net_10153;
wire net_3119;
wire net_1231;
wire net_5841;
wire net_19009;
wire net_6205;
wire net_815;
wire net_7875;
wire net_18951;
wire net_11304;
wire net_15049;
wire net_18022;
wire x186;
wire net_6514;
wire net_7897;
wire net_7670;
wire net_5632;
wire net_10279;
wire net_586;
wire net_10845;
wire net_1347;
wire net_1091;
wire net_15926;
wire net_13145;
wire net_16724;
wire net_18112;
wire net_3745;
wire net_11713;
wire net_9879;
wire net_16030;
wire net_3708;
wire net_5830;
wire net_5227;
wire net_7536;
wire net_14259;
wire net_7042;
wire net_6073;
wire net_7478;
wire net_16302;
wire net_16202;
wire net_2556;
wire net_8599;
wire net_16271;
wire net_3519;
wire net_2740;
wire net_14756;
wire net_7294;
wire net_672;
wire net_18548;
wire net_15015;
wire net_8834;
wire net_5212;
wire net_16938;
wire net_16914;
wire net_2027;
wire net_13761;
wire net_11680;
wire net_7021;
wire net_3610;
wire net_8963;
wire net_5784;
wire net_1953;
wire net_15177;
wire net_17630;
wire net_14295;
wire net_3925;
wire net_3847;
wire net_4473;
wire net_8230;
wire net_4582;
wire net_18339;
wire net_4547;
wire net_14205;
wire net_7819;
wire net_14455;
wire net_8954;
wire net_15154;
wire net_18837;
wire net_10136;
wire net_16776;
wire net_4640;
wire net_17520;
wire net_10926;
wire net_11602;
wire x13482;
wire net_7071;
wire net_7982;
wire net_13264;
wire net_802;
wire net_16610;
wire net_12194;
wire net_12930;
wire net_4997;
wire net_14359;
wire net_9230;
wire net_6620;
wire net_17817;
wire net_17784;
wire net_4824;
wire net_15181;
wire net_7049;
wire net_14189;
wire net_13404;
wire net_1636;
wire net_7568;
wire net_9714;
wire net_16293;
wire net_3257;
wire net_4458;
wire net_10899;
wire net_10344;
wire net_10270;
wire net_16777;
wire net_1334;
wire net_18374;
wire net_10782;
wire net_757;
wire net_206;
wire net_10087;
wire net_10894;
wire net_15430;
wire net_14134;
wire net_235;
wire net_13121;
wire net_14970;
wire net_11695;
wire net_12223;
wire net_2961;
wire net_18775;
wire net_5108;
wire net_7652;
wire net_5631;
wire net_3644;
wire net_16333;
wire net_12273;
wire net_3081;
wire net_12927;
wire net_11279;
wire net_10283;
wire net_4879;
wire net_6144;
wire net_17842;
wire net_14570;
wire net_2630;
wire net_1985;
wire net_2340;
wire net_14421;
wire net_14883;
wire net_2275;
wire net_10752;
wire net_3976;
wire net_9619;
wire net_10939;
wire net_13128;
wire net_841;
wire net_10803;
wire net_1750;
wire net_6411;
wire net_3346;
wire x13750;
wire net_8269;
wire net_528;
wire net_335;
wire net_4878;
wire net_15778;
wire net_3464;
wire net_9132;
wire net_181;
wire net_9661;
wire net_6784;
wire net_15796;
wire net_12214;
wire net_3333;
wire net_11556;
wire net_6011;
wire net_10631;
wire net_9014;
wire net_13530;
wire net_6177;
wire net_3649;
wire net_2539;
wire net_18055;
wire net_17555;
wire net_6216;
wire net_386;
wire net_12680;
wire net_6150;
wire net_10051;
wire net_1790;
wire net_8166;
wire net_4103;
wire net_11221;
wire net_6130;
wire net_15719;
wire net_10583;
wire net_12718;
wire net_7573;
wire net_1709;
wire net_10981;
wire net_10080;
wire net_17294;
wire net_9698;
wire net_5707;
wire net_18404;
wire net_13622;
wire net_175;
wire net_12650;
wire net_1850;
wire net_4429;
wire net_6365;
wire net_1992;
wire net_15606;
wire net_17377;
wire net_12346;
wire net_897;
wire net_7384;
wire net_11362;
wire net_2853;
wire net_10578;
wire net_2705;
wire net_5164;
wire net_615;
wire net_6712;
wire net_18104;
wire net_441;
wire net_16338;
wire net_14224;
wire net_17564;
wire net_17279;
wire net_6032;
wire net_17627;
wire net_2663;
wire net_17949;
wire net_728;
wire net_1276;
wire net_5473;
wire net_7774;
wire net_14905;
wire net_170;
wire net_17353;
wire net_15138;
wire net_16495;
wire net_5305;
wire net_10741;
wire net_17299;
wire net_17050;
wire net_16986;
wire net_14661;
wire net_3321;
wire net_15836;
wire net_15342;
wire net_15631;
wire net_13764;
wire net_708;
wire net_7685;
wire net_16667;
wire net_3216;
wire net_171;
wire net_9796;
wire net_16631;
wire net_15134;
wire net_10013;
wire net_6563;
wire net_10528;
wire net_18289;
wire net_604;
wire net_14578;
wire net_17322;
wire net_15465;
wire net_16507;
wire net_12385;
wire net_483;
wire net_15439;
wire net_16519;
wire net_1149;
wire net_9937;
wire net_8097;
wire net_15507;
wire net_16283;
wire net_16025;
wire net_15318;
wire net_2131;
wire net_6681;
wire net_16568;
wire x729;
wire net_5651;
wire net_13461;
wire net_12845;
wire net_18484;
wire net_15981;
wire net_7153;
wire net_13632;
wire net_11369;
wire net_2228;
wire net_12357;
wire net_786;
wire net_5141;
wire net_11801;
wire net_11564;
wire net_8998;
wire net_17308;
wire net_9470;
wire net_17896;
wire net_9892;
wire net_9080;
wire net_8461;
wire net_3577;
wire net_10137;
wire net_1815;
wire net_3840;
wire net_4361;
wire net_15458;
wire net_6145;
wire net_3782;
wire net_13250;
wire net_877;
wire net_14680;
wire net_2799;
wire net_6868;
wire net_6834;
wire net_8092;
wire net_3734;
wire net_14135;
wire net_14524;
wire net_8021;
wire net_15714;
wire net_9654;
wire net_11570;
wire net_11232;
wire net_4066;
wire net_13296;
wire net_6257;
wire net_14869;
wire net_8026;
wire net_3284;
wire net_1474;
wire net_4297;
wire net_18675;
wire net_15482;
wire net_12088;
wire net_2784;
wire net_17108;
wire net_15642;
wire net_13843;
wire net_8753;
wire net_675;
wire net_8355;
wire net_2867;
wire net_3472;
wire net_9120;
wire net_10700;
wire net_7578;
wire x3904;
wire net_1768;
wire net_16010;
wire net_12950;
wire net_7677;
wire net_304;
wire net_17968;
wire net_16427;
wire net_9791;
wire net_7326;
wire net_14967;
wire net_4347;
wire net_10551;
wire net_7731;
wire net_15431;
wire net_18660;
wire net_12731;
wire net_15517;
wire net_1316;
wire net_6845;
wire net_6545;
wire net_17311;
wire net_792;
wire net_15744;
wire net_13848;
wire net_6223;
wire net_13782;
wire net_8842;
wire net_2203;
wire net_4430;
wire net_13415;
wire net_5373;
wire net_5678;
wire net_18635;
wire net_18242;
wire net_219;
wire net_3609;
wire net_18125;
wire net_9976;
wire net_2476;
wire net_15791;
wire net_13798;
wire net_913;
wire net_4518;
wire net_5378;
wire net_5338;
wire net_14938;
wire net_13591;
wire net_15423;
wire net_4330;
wire net_7756;
wire net_4019;
wire net_15037;
wire net_4152;
wire net_10832;
wire net_360;
wire net_13561;
wire net_7017;
wire net_14832;
wire net_2324;
wire net_18925;
wire net_11688;
wire net_16961;
wire net_4805;
wire net_13259;
wire net_3316;
wire net_10162;
wire net_3032;
wire net_9507;
wire net_17484;
wire net_1373;
wire net_1352;
wire net_2885;
wire net_16605;
wire net_10735;
wire net_4696;
wire net_17127;
wire net_8814;
wire net_17087;
wire net_1187;
wire net_17079;
wire net_7408;
wire net_4988;
wire net_3206;
wire net_17163;
wire net_2858;
wire net_18696;
wire net_15470;
wire net_14806;
wire net_14703;
wire net_15004;
wire net_5569;
wire net_12234;
wire net_12047;
wire net_1442;
wire net_18410;
wire net_16400;
wire net_10042;
wire net_11544;
wire net_15188;
wire net_16968;
wire net_17411;
wire net_12298;
wire net_1894;
wire net_9645;
wire net_10694;
wire net_2431;
wire net_8213;
wire net_633;
wire net_5750;
wire net_10115;
wire net_1914;
wire x12780;
wire net_15996;
wire net_14944;
wire net_2408;
wire net_9904;
wire net_6627;
wire net_5943;
wire net_6974;
wire net_15022;
wire net_14669;
wire net_15540;
wire net_1457;
wire net_2741;
wire net_7010;
wire net_18982;
wire net_5414;
wire net_14876;
wire net_4011;
wire net_17721;
wire net_1436;
wire net_9199;
wire net_4338;
wire net_10054;
wire net_10725;
wire net_3392;
wire net_9571;
wire net_2551;
wire net_11572;
wire net_12547;
wire net_14348;
wire net_6323;
wire net_2891;
wire net_14314;
wire net_8928;
wire net_11261;
wire net_15269;
wire net_18672;
wire net_2401;
wire net_14502;
wire x1829;
wire net_15530;
wire net_1305;
wire net_17735;
wire net_16482;
wire x831;
wire net_14493;
wire net_1387;
wire net_1581;
wire net_11808;
wire net_4468;
wire net_2413;
wire net_7786;
wire net_14462;
wire net_2792;
wire net_345;
wire net_2965;
wire net_2128;
wire net_16722;
wire net_9990;
wire net_17438;
wire net_11891;
wire net_5302;
wire net_11489;
wire net_9344;
wire net_5080;
wire net_11140;
wire net_17219;
wire net_13584;
wire net_2461;
wire net_14654;
wire net_1766;
wire net_2582;
wire net_8974;
wire net_7898;
wire net_10419;
wire net_3872;
wire net_4956;
wire net_17098;
wire net_11867;
wire net_19027;
wire net_9407;
wire net_4447;
wire net_10357;
wire net_15826;
wire net_10226;
wire net_13933;
wire net_9235;
wire net_8990;
wire net_14166;
wire net_8794;
wire net_9834;
wire net_12667;
wire net_13536;
wire net_13443;
wire net_17155;
wire net_10387;
wire net_1759;
wire net_12996;
wire net_15308;
wire net_12752;
wire net_3764;
wire net_12964;
wire net_18395;
wire net_11636;
wire net_2541;
wire net_12310;
wire net_3689;
wire net_12635;
wire net_533;
wire net_7436;
wire net_911;
wire net_7775;
wire net_12017;
wire net_10047;
wire net_9608;
wire net_6637;
wire net_9015;
wire net_7053;
wire net_5570;
wire net_15463;
wire net_11745;
wire net_9457;
wire net_13709;
wire net_7962;
wire net_17981;
wire net_6485;
wire net_5312;
wire net_5861;
wire net_18182;
wire net_1443;
wire net_16699;
wire net_11888;
wire net_8691;
wire net_18815;
wire net_16498;
wire net_2840;
wire net_16929;
wire net_14721;
wire net_3463;
wire net_4005;
wire net_6008;
wire net_17910;
wire net_16763;
wire net_11883;
wire net_3199;
wire net_8001;
wire net_3597;
wire net_5671;
wire net_15602;
wire net_16422;
wire net_269;
wire net_5043;
wire net_3193;
wire net_3131;
wire net_10107;
wire net_12171;
wire net_3179;
wire net_1945;
wire net_10064;
wire net_7207;
wire net_10858;
wire net_4073;
wire net_5159;
wire net_1833;
wire x4214;
wire net_8496;
wire net_2831;
wire net_3029;
wire net_18296;
wire net_9622;
wire net_7818;
wire net_5725;
wire net_12779;
wire net_8252;
wire net_18688;
wire net_6523;
wire net_17182;
wire net_5064;
wire net_6024;
wire net_17876;
wire net_11780;
wire net_12154;
wire net_15755;
wire net_8172;
wire net_7912;
wire net_16408;
wire net_5380;
wire net_10173;
wire net_8519;
wire net_5648;
wire net_14246;
wire net_18006;
wire net_11152;
wire net_16147;
wire net_11251;
wire net_10644;
wire net_3980;
wire net_10566;
wire net_1481;
wire net_10392;
wire net_7922;
wire net_16875;
wire x808;
wire net_700;
wire net_5000;
wire net_11433;
wire net_9947;
wire net_11043;
wire net_6043;
wire net_18300;
wire net_5216;
wire net_15195;
wire net_18681;
wire net_11819;
wire net_1673;
wire net_11941;
wire net_3480;
wire net_6715;
wire net_8933;
wire net_4135;
wire net_6982;
wire net_2945;
wire net_17826;
wire net_16682;
wire net_12855;
wire net_3665;
wire net_717;
wire net_544;
wire net_15587;
wire net_12305;
wire net_10505;
wire net_15328;
wire net_8201;
wire net_9659;
wire net_18251;
wire net_3402;
wire net_2223;
wire net_6957;
wire net_8008;
wire net_2673;
wire net_3500;
wire net_6164;
wire net_9358;
wire net_5903;
wire x677;
wire net_17706;
wire net_1245;
wire net_3660;
wire net_5806;
wire net_18632;
wire net_870;
wire net_7135;
wire net_7176;
wire net_7521;
wire net_10819;
wire net_7941;
wire net_13642;
wire net_12012;
wire net_14581;
wire net_6286;
wire net_17855;
wire net_12874;
wire net_12668;
wire net_11645;
wire net_5127;
wire net_17031;
wire net_14155;
wire net_10922;
wire net_7362;
wire net_14084;
wire net_16649;
wire net_19015;
wire net_2920;
wire net_1591;
wire net_7695;
wire net_1747;
wire net_650;
wire x1667;
wire net_15080;
wire net_9761;
wire net_597;
wire net_17852;
wire net_14065;
wire net_17321;
wire x3983;
wire net_15767;
wire net_5984;
wire net_10482;
wire net_8272;
wire x291;
wire net_15109;
wire net_14281;
wire net_6336;
wire x508;
wire net_12481;
wire net_8889;
wire net_10853;
wire net_18161;
wire net_19026;
wire net_603;
wire net_4913;
wire net_642;
wire net_16314;
wire net_9806;
wire net_2699;
wire net_1158;
wire net_6989;
wire net_11496;
wire net_8006;
wire net_11082;
wire net_10775;
wire net_11530;
wire net_13964;
wire net_470;
wire net_2702;
wire net_430;
wire net_2834;
wire net_11659;
wire net_15255;
wire net_17442;
wire net_17346;
wire net_15903;
wire x4323;
wire net_3129;
wire x13252;
wire net_18526;
wire net_8568;
wire net_12353;
wire net_18797;
wire net_11771;
wire net_1063;
wire net_4218;
wire net_14644;
wire net_12571;
wire net_18546;
wire net_9127;
wire net_7297;
wire net_13577;
wire net_15089;
wire net_17763;
wire net_1504;
wire net_475;
wire net_6737;
wire net_9432;
wire net_7216;
wire net_14272;
wire net_11137;
wire net_14024;
wire net_13768;
wire net_6903;
wire net_2470;
wire net_11474;
wire net_1568;
wire net_14288;
wire x2856;
wire net_6756;
wire net_1526;
wire net_13860;
wire net_1884;
wire net_12341;
wire net_3919;
wire net_16920;
wire net_2646;
wire net_3936;
wire net_4364;
wire net_13198;
wire net_6645;
wire net_17538;
wire net_1360;
wire net_6344;
wire net_3364;
wire net_5316;
wire net_14420;
wire net_1364;
wire net_6003;
wire net_5050;
wire net_14727;
wire net_17550;
wire net_827;
wire net_549;
wire net_10192;
wire net_11050;
wire net_4563;
wire net_2337;
wire net_14928;
wire net_6945;
wire net_1369;
wire net_6900;
wire net_11068;
wire net_4695;
wire net_8622;
wire net_1013;
wire net_16865;
wire net_1530;
wire net_16345;
wire net_16809;
wire net_13869;
wire net_3075;
wire net_842;
wire net_11783;
wire net_2336;
wire net_1705;
wire net_14977;
wire net_6571;
wire net_9500;
wire x886;
wire net_11215;
wire net_8951;
wire net_6560;
wire net_10325;
wire net_8199;
wire net_3739;
wire net_8455;
wire net_492;
wire net_11392;
wire net_3678;
wire net_7234;
wire net_8797;
wire net_2639;
wire net_8071;
wire net_16085;
wire net_13370;
wire net_16702;
wire net_3695;
wire net_5450;
wire net_1327;
wire net_17650;
wire net_4968;
wire net_15337;
wire net_12734;
wire net_2248;
wire net_4971;
wire net_11532;
wire net_3866;
wire net_6772;
wire net_13473;
wire net_7787;
wire net_13223;
wire net_14548;
wire net_12024;
wire net_12920;
wire net_4300;
wire net_9578;
wire net_4776;
wire net_17676;
wire net_10477;
wire net_15167;
wire net_13820;
wire net_2868;
wire net_6083;
wire net_16037;
wire net_15074;
wire net_8295;
wire net_2946;
wire net_11373;
wire net_1284;
wire net_4397;
wire x2981;
wire net_13977;
wire net_13732;
wire net_13095;
wire net_6671;
wire net_16376;
wire net_3929;
wire net_16321;
wire net_9942;
wire net_13888;
wire net_7567;
wire net_15536;
wire net_18530;
wire net_17422;
wire net_16477;
wire net_2066;
wire net_18439;
wire net_13925;
wire net_9310;
wire net_7415;
wire net_8109;
wire net_1146;
wire net_11679;
wire net_4612;
wire net_15815;
wire net_4519;
wire net_17671;
wire net_18097;
wire net_16905;
wire net_8584;
wire net_16739;
wire net_13881;
wire net_17239;
wire net_16015;
wire net_9897;
wire net_18933;
wire net_5495;
wire net_13071;
wire net_9511;
wire net_8284;
wire net_2762;
wire net_17525;
wire net_11828;
wire net_6439;
wire net_6247;
wire net_14569;
wire net_6424;
wire net_4619;
wire net_6377;
wire net_10161;
wire net_2089;
wire net_6352;
wire net_12429;
wire net_3797;
wire net_15391;
wire net_9718;
wire net_3535;
wire net_12248;
wire net_1195;
wire net_18174;
wire net_17884;
wire net_16821;
wire net_2502;
wire net_1396;
wire net_16919;
wire net_4069;
wire x13921;
wire net_7225;
wire x4733;
wire net_2737;
wire net_6397;
wire net_5126;
wire net_18515;
wire net_18408;
wire net_14828;
wire net_12108;
wire net_2481;
wire net_4539;
wire net_15698;
wire net_15094;
wire net_10624;
wire net_8104;
wire net_14210;
wire net_17134;
wire x2230;
wire net_2617;
wire net_1060;
wire net_12699;
wire net_4846;
wire x494;
wire net_12101;
wire net_1715;
wire net_15961;
wire net_9913;
wire net_14842;
wire net_7583;
wire net_9234;
wire net_15221;
wire net_14557;
wire net_6577;
wire net_1216;
wire net_4599;
wire net_14583;
wire net_2815;
wire net_15040;
wire net_3785;
wire net_18994;
wire net_11240;
wire net_1271;
wire net_1086;
wire net_18465;
wire net_9593;
wire net_10978;
wire net_13453;
wire net_1197;
wire net_7613;
wire net_5744;
wire net_5858;
wire net_11752;
wire net_18018;
wire net_576;
wire net_8932;
wire net_1654;
wire x794;
wire net_8438;
wire net_3005;
wire net_11183;
wire net_12902;
wire net_10679;
wire net_11272;
wire net_725;
wire net_3931;
wire net_17591;
wire net_18369;
wire net_6183;
wire net_14766;
wire net_894;
wire net_16219;
wire net_13914;
wire net_10545;
wire x13712;
wire net_17718;
wire net_18496;
wire net_1423;
wire net_13012;
wire net_2902;
wire net_1871;
wire net_517;
wire net_628;
wire net_18030;
wire net_3494;
wire net_6600;
wire net_12123;
wire net_10377;
wire net_14018;
wire net_10204;
wire net_9555;
wire net_9036;
wire net_17482;
wire net_17691;
wire net_6406;
wire net_10322;
wire net_1289;
wire x13018;
wire net_3138;
wire net_14858;
wire net_11982;
wire net_15786;
wire net_13377;
wire net_12867;
wire net_6922;
wire net_17061;
wire net_11162;
wire net_5895;
wire net_12446;
wire net_5876;
wire x13100;
wire net_2723;
wire net_17365;
wire net_15144;
wire net_5157;
wire net_13504;
wire net_2552;
wire net_3229;
wire net_1001;
wire net_13778;
wire net_781;
wire net_3765;
wire net_8479;
wire net_15323;
wire net_13063;
wire net_5241;
wire net_7506;
wire net_5967;
wire x13396;
wire net_6818;
wire net_16677;
wire net_13188;
wire net_16353;
wire net_185;
wire net_7357;
wire net_17195;
wire net_16194;
wire net_14687;
wire net_16540;
wire net_4321;
wire net_4631;
wire net_18452;
wire net_1015;
wire net_2980;
wire net_14685;
wire net_16717;
wire net_9863;
wire net_9772;
wire net_11964;
wire net_5794;
wire net_14748;
wire net_7766;
wire net_17489;
wire net_11759;
wire net_6856;
wire net_15660;
wire net_2146;
wire net_405;
wire net_11927;
wire net_1111;
wire net_11614;
wire net_2651;
wire net_4281;
wire net_8259;
wire net_3971;
wire net_16841;
wire net_16224;
wire net_3155;
wire net_7969;
wire net_831;
wire net_4728;
wire net_5442;
wire net_451;
wire net_1234;
wire net_750;
wire net_12558;
wire net_7835;
wire net_9746;
wire net_16411;
wire net_13027;
wire net_12797;
wire net_7274;
wire net_17866;
wire net_17274;
wire net_14641;
wire net_11459;
wire net_8571;
wire net_5915;
wire net_18738;
wire net_5184;
wire net_17401;
wire x2133;
wire net_16189;
wire x1500;
wire net_5788;
wire net_11920;
wire net_8472;
wire net_773;
wire net_4759;
wire net_11770;
wire net_9590;
wire net_16653;
wire net_11796;
wire net_11622;
wire net_8537;
wire net_12098;
wire net_15976;
wire net_3727;
wire net_15887;
wire net_13986;
wire net_6766;
wire net_13269;
wire net_6355;
wire net_5052;
wire net_14400;
wire net_9997;
wire net_8305;
wire net_14091;
wire net_4205;
wire net_834;
wire net_10298;
wire net_694;
wire net_13615;
wire net_13556;
wire net_18528;
wire net_13794;
wire net_5925;
wire net_9950;
wire net_7609;
wire net_8778;
wire net_8946;
wire net_8409;
wire net_1570;
wire net_13385;
wire net_4645;
wire net_11100;
wire net_17415;
wire net_12204;
wire net_9499;
wire net_11228;
wire net_7320;
wire net_15811;
wire net_8779;
wire net_252;
wire net_10497;
wire net_7693;
wire net_14897;
wire net_2399;
wire net_16325;
wire net_14508;
wire net_901;
wire net_6267;
wire net_7846;
wire net_3425;
wire net_16780;
wire net_410;
wire net_8134;
wire net_4243;
wire net_14940;
wire net_10539;
wire net_9136;
wire net_6798;
wire net_6607;
wire net_12470;
wire net_18956;
wire net_7886;
wire net_17473;
wire net_2603;
wire net_5910;
wire net_7824;
wire net_1132;
wire net_14144;
wire net_5880;
wire net_10351;
wire net_2442;
wire net_3026;
wire net_7743;
wire net_13749;
wire net_12317;
wire net_9410;
wire net_5760;
wire net_18869;
wire net_5923;
wire net_2356;
wire net_3288;
wire net_971;
wire net_8194;
wire net_11734;
wire net_2184;
wire net_18278;
wire net_11824;
wire net_554;
wire net_16894;
wire net_14544;
wire net_13625;
wire net_18765;
wire net_4653;
wire net_14232;
wire net_11187;
wire net_8704;
wire net_3740;
wire net_15278;
wire net_14221;
wire net_8317;
wire net_6306;
wire net_584;
wire net_13753;
wire net_10446;
wire net_12656;
wire net_2411;
wire net_13104;
wire net_11511;
wire net_165;
wire net_9226;
wire net_16055;
wire net_14794;
wire net_18585;
wire net_3438;
wire net_3824;
wire net_8789;
wire net_4440;
wire net_8576;
wire net_18847;
wire net_13612;
wire net_10170;
wire net_16215;
wire net_12970;
wire net_3823;
wire net_9886;
wire net_17888;
wire net_8600;
wire net_18970;
wire net_16832;
wire net_17795;
wire net_9365;
wire net_13573;
wire net_3859;
wire net_8044;
wire net_15350;
wire net_7885;
wire net_3803;
wire net_17664;
wire net_8607;
wire net_11284;
wire net_16099;
wire net_15395;
wire net_14338;
wire net_14592;
wire net_8880;
wire net_8592;
wire net_7707;
wire net_3334;
wire net_6789;
wire net_3224;
wire net_1719;
wire net_17740;
wire net_15613;
wire net_15854;
wire net_16068;
wire net_5715;
wire net_11562;
wire net_15739;
wire net_11464;
wire net_15426;
wire net_8786;
wire net_17917;
wire net_14448;
wire net_8034;
wire net_11598;
wire net_2440;
wire net_9386;
wire net_18995;
wire net_16077;
wire x13353;
wire net_6809;
wire net_14043;
wire net_12800;
wire net_1379;
wire x13779;
wire net_1322;
wire net_14437;
wire net_9538;
wire net_8526;
wire x13520;
wire net_12143;
wire net_10373;
wire net_1301;
wire net_12066;
wire net_14258;
wire net_12487;
wire net_8749;
wire x13698;
wire net_7596;
wire net_12756;
wire net_7247;
wire net_6932;
wire net_7116;
wire net_16575;
wire net_17456;
wire net_426;
wire net_5203;
wire net_16298;
wire net_6095;
wire net_14511;
wire net_414;
wire net_7793;
wire net_17611;
wire net_1048;
wire net_18249;
wire net_3048;
wire net_799;
wire net_5102;
wire net_5576;
wire net_18057;
wire net_15367;
wire net_5737;
wire net_12588;
wire net_2014;
wire x863;
wire net_16884;
wire net_16278;
wire net_6747;
wire net_13487;
wire net_5999;
wire net_9845;
wire net_16952;
wire net_4742;
wire net_2454;
wire net_8917;
wire net_8716;
wire net_4761;
wire net_14709;
wire net_17547;
wire net_18151;
wire net_7616;
wire net_15701;
wire net_16582;
wire net_6016;
wire net_18498;
wire net_17603;
wire net_10140;
wire net_15972;
wire net_12621;
wire net_247;
wire net_14630;
wire x13576;
wire net_3413;
wire net_14430;
wire net_9742;
wire net_8619;
wire net_12627;
wire net_1934;
wire net_14180;
wire net_13740;
wire net_12513;
wire net_6235;
wire net_11327;
wire net_1848;
wire x919;
wire net_639;
wire net_4724;
wire net_9583;
wire net_18363;
wire net_12309;
wire net_5697;
wire net_1238;
wire net_14923;
wire net_13697;
wire net_14074;
wire net_7599;
wire net_9483;
wire net_1033;
wire net_10604;
wire net_5560;
wire net_12458;
wire net_11333;
wire net_8333;
wire net_13149;
wire net_15163;
wire net_12005;
wire net_12302;
wire net_3107;
wire net_7069;
wire net_1686;
wire net_11860;
wire net_11481;
wire net_10686;
wire net_10263;
wire x3207;
wire net_367;
wire net_3303;
wire net_17861;
wire net_17747;
wire net_6296;
wire net_10061;
wire net_1842;
wire net_9849;
wire net_13037;
wire net_8774;
wire net_3957;
wire net_1180;
wire net_8561;
wire net_1627;
wire net_10235;
wire net_5869;
wire net_2002;
wire net_1069;
wire net_2022;
wire net_9932;
wire net_12014;
wire net_5406;
wire net_18591;
wire net_2385;
wire net_3431;
wire net_17118;
wire net_5829;
wire net_3565;
wire net_7009;
wire net_1416;
wire net_7656;
wire net_13484;
wire net_18167;
wire net_6065;
wire net_2433;
wire net_15111;
wire net_6726;
wire net_4029;
wire net_1601;
wire net_6614;
wire net_4087;
wire net_4255;
wire net_9854;
wire net_17659;
wire net_13437;
wire net_8866;
wire net_348;
wire net_7398;
wire net_9667;
wire net_626;
wire net_10796;
wire net_15260;
wire net_5068;
wire net_16116;
wire net_11257;
wire net_1809;
wire net_686;
wire net_17904;
wire net_1615;
wire net_16521;
wire net_17266;
wire net_14037;
wire net_17192;
wire net_7859;
wire net_17495;
wire net_4578;
wire net_2112;
wire net_5072;
wire net_14505;
wire net_1828;
wire net_16063;
wire net_1466;
wire net_5320;
wire net_10438;
wire net_16182;
wire net_11268;
wire net_157;
wire net_17074;
wire net_6695;
wire net_9006;
wire net_7759;
wire net_18139;
wire net_1205;
wire net_11627;
wire net_8154;
wire net_6978;
wire net_466;
wire net_9612;
wire net_1179;
wire net_18232;
wire net_15844;
wire net_15231;
wire net_18720;
wire net_7833;
wire net_13057;
wire net_16709;
wire net_11021;
wire net_16289;
wire net_1610;
wire net_3569;
wire net_6814;
wire net_13236;
wire net_4246;
wire net_8893;
wire net_4020;
wire net_16870;
wire net_8389;
wire net_4453;
wire net_17282;
wire net_16467;
wire net_15593;
wire net_11018;
wire net_7118;
wire net_644;
wire net_13495;
wire net_12111;
wire net_12063;
wire net_852;
wire net_11917;
wire net_11035;
wire net_15118;
wire net_14771;
wire net_7391;
wire net_8904;
wire net_8416;
wire net_8382;
wire net_11404;
wire net_18706;
wire net_14690;
wire net_14284;
wire net_10128;
wire net_8685;
wire net_11492;
wire net_9491;
wire net_8555;
wire net_11410;
wire net_5871;
wire net_14061;
wire net_15243;
wire net_1693;
wire net_10707;
wire net_8853;
wire net_3779;
wire net_4252;
wire net_2068;
wire net_17880;
wire net_14659;
wire net_3705;
wire net_5907;
wire net_11821;
wire net_16673;
wire x703;
wire net_5930;
wire net_6371;
wire net_8939;
wire net_17584;
wire net_15692;
wire net_314;
wire net_5395;
wire net_17637;
wire net_15301;
wire net_18615;
wire net_11381;
wire net_9765;
wire net_18623;
wire net_12033;
wire net_14964;
wire net_8442;
wire net_4669;
wire x13457;
wire net_13791;
wire net_5460;
wire net_12479;
wire net_4286;
wire net_9872;
wire net_3484;
wire net_16518;
wire net_945;
wire net_6532;
wire net_4380;
wire net_6971;
wire net_12266;
wire net_2101;
wire net_7738;
wire net_6863;
wire net_18572;
wire net_11451;
wire net_8875;
wire net_8376;
wire net_15246;
wire net_6582;
wire net_5800;
wire net_5601;
wire net_15312;
wire net_13426;
wire net_16851;
wire net_12251;
wire net_8808;
wire net_6340;
wire net_13256;
wire net_10516;
wire net_18823;
wire net_9099;
wire net_5174;
wire net_11343;
wire net_8943;
wire net_1784;
wire net_1296;
wire net_17253;
wire net_15738;
wire net_16823;
wire net_13081;
wire net_4326;
wire net_10245;
wire net_7159;
wire net_10762;
wire net_9735;
wire net_2424;
wire net_1968;
wire net_15364;
wire net_10746;
wire net_10407;
wire net_12291;
wire net_4488;
wire net_5092;
wire net_5295;
wire net_18534;
wire net_7713;
wire net_2507;
wire net_17024;
wire net_16791;
wire net_9633;
wire net_17335;
wire net_13908;
wire net_2685;
wire net_8340;
wire net_14264;
wire net_2898;
wire net_6197;
wire net_1391;
wire net_9334;
wire net_14933;
wire net_9926;
wire net_5132;
wire net_18203;
wire x12991;
wire net_10304;
wire net_17235;
wire net_14847;
wire net_1772;
wire net_14552;
wire net_3529;
wire net_6128;
wire net_5437;
wire net_2498;
wire net_381;
wire net_9144;
wire net_6574;
wire net_6889;
wire net_10710;
wire net_15891;
wire net_3783;
wire net_1857;
wire net_7445;
wire net_11586;
wire net_11010;
wire net_12059;
wire net_6109;
wire net_15554;
wire net_14414;
wire net_9883;
wire net_17993;
wire net_16751;
wire net_1557;
wire net_6843;
wire net_1514;
wire net_3852;
wire net_7668;
wire net_13072;
wire net_6825;
wire net_13874;
wire net_3092;
wire net_14407;
wire net_9209;
wire net_8802;
wire net_6995;
wire net_13240;
wire net_12241;
wire net_500;
wire net_5357;
wire net_1906;
wire net_17687;
wire net_9094;
wire net_8056;
wire net_5660;
wire net_15410;
wire net_11967;
wire net_14197;
wire net_10911;
wire net_14120;
wire net_17822;
wire net_14717;
wire net_10130;
wire net_11974;
wire net_16992;
wire net_4401;
wire net_18355;
wire net_15271;
wire net_3632;
wire net_2189;
wire net_2057;
wire net_1124;
wire net_13945;
wire net_7645;
wire net_16816;
wire net_13737;
wire net_5960;
wire net_5615;
wire net_143;
wire net_12434;
wire net_190;
wire net_4964;
wire net_1447;
wire net_1929;
wire net_9423;
wire net_3493;
wire net_2061;
wire net_13466;
wire net_5288;
wire net_15878;
wire net_13956;
wire net_14030;
wire net_13910;
wire net_13727;
wire net_14780;
wire net_13710;
wire net_1895;
wire net_5360;
wire net_509;
wire net_14983;
wire net_4975;
wire net_16157;
wire net_9983;
wire net_211;
wire net_16248;
wire net_13430;
wire net_10079;
wire net_6752;
wire net_14564;
wire net_18001;
wire net_5771;
wire net_13541;
wire net_3941;
wire net_6630;
wire net_12604;
wire net_17359;
wire net_8645;
wire net_2233;
wire net_2033;
wire net_18061;
wire net_12726;
wire net_12091;
wire net_8487;
wire net_15710;
wire net_2123;
wire net_10811;
wire net_12784;
wire net_12360;
wire net_9049;
wire net_5970;
wire net_16554;
wire net_2532;
wire x13004;
wire net_18468;
wire net_12785;
wire net_13851;
wire net_11112;
wire net_1864;
wire net_15441;
wire net_14917;
wire net_11725;
wire net_6156;
wire net_12840;
wire net_2518;
wire net_14604;
wire net_6950;
wire net_10663;
wire net_4062;
wire x926;
wire net_17014;
wire net_12284;
wire net_14353;
wire net_7953;
wire net_1646;
wire net_4115;
wire net_11437;
wire net_2776;
wire net_18433;
wire net_3389;
wire net_12938;
wire net_1562;
wire net_16743;
wire net_15225;
wire net_2522;
wire net_4178;
wire net_7267;
wire net_8671;
wire net_17928;
wire net_13878;
wire net_12987;
wire net_1524;
wire net_16398;
wire net_18385;
wire net_10022;
wire net_9396;
wire net_17943;
wire net_15686;
wire net_12531;
wire net_9785;
wire net_11670;
wire net_15864;
wire net_16572;
wire net_6461;
wire net_2511;
wire net_2626;
wire net_2115;
wire net_4110;
wire net_4317;
wire net_2299;
wire net_9307;
wire net_10612;
wire net_16049;
wire net_7123;
wire net_17837;
wire net_1405;
wire net_7726;
wire net_10072;
wire net_17902;
wire net_13518;
wire net_10881;
wire net_6555;
wire net_15102;
wire net_716;
wire net_5147;
wire net_13273;
wire net_13200;
wire net_10489;
wire net_11445;
wire net_1269;
wire net_16846;
wire net_13757;
wire net_8630;
wire net_3715;
wire net_3533;
wire net_5400;
wire net_11805;
wire net_12406;
wire net_4293;
wire net_9176;
wire net_666;
wire net_13776;
wire net_4809;
wire net_11308;
wire net_18305;
wire net_12706;
wire net_12184;
wire net_6212;
wire net_9702;
wire net_15125;
wire net_3946;
wire net_10596;
wire net_5522;
wire net_6319;
wire net_7636;
wire net_9024;
wire net_9824;
wire net_1657;
wire net_6063;
wire net_3084;
wire net_10689;
wire net_10863;
wire net_19010;
wire net_18894;
wire net_18477;
wire net_17380;
wire net_9859;
wire net_3994;
wire net_18790;
wire net_11764;
wire net_14213;
wire net_13645;
wire net_1976;
wire net_8510;
wire net_3169;
wire net_14734;
wire net_5647;
wire net_3792;
wire x1244;
wire net_2758;
wire net_9972;
wire net_1826;
wire net_18327;
wire net_14634;
wire net_16531;
wire net_4609;
wire net_10337;
wire net_16860;
wire net_16160;
wire net_2142;
wire net_11841;
wire net_15335;
wire net_7332;
wire net_920;
wire net_3009;
wire net_12980;
wire net_5596;
wire net_15653;
wire net_4226;
wire net_820;
wire net_7137;
wire net_18656;
wire net_11249;
wire net_16530;
wire net_15765;
wire x697;
wire net_18901;
wire net_13447;
wire net_6137;
wire net_13465;
wire net_5959;
wire net_9681;
wire net_566;
wire net_5063;
wire net_7519;
wire net_9768;
wire net_13173;
wire net_13811;
wire net_4735;
wire net_17771;
wire net_18788;
wire net_17696;
wire net_2108;
wire net_2529;
wire net_19038;
wire net_6044;
wire net_4685;
wire net_4732;
wire net_9751;
wire net_8390;
wire x1977;
wire net_5979;
wire net_7551;
wire net_11810;
wire net_18985;
wire net_18024;
wire net_14279;
wire net_4235;
wire net_15570;
wire net_14117;
wire net_11871;
wire net_14990;
wire net_13379;
wire net_9452;
wire net_4117;
wire net_1357;
wire net_15875;
wire net_13990;
wire net_3637;
wire net_5554;
wire net_18564;
wire net_17188;
wire net_14476;
wire net_8668;
wire net_18966;
wire net_4604;
wire net_7489;
wire net_6558;
wire net_12598;
wire net_419;
wire net_12463;
wire net_16974;
wire net_5658;
wire net_936;
wire net_15400;
wire net_9259;
wire net_8066;
wire net_7808;
wire net_17006;
wire x13833;
wire net_819;
wire net_10969;
wire net_11954;
wire net_8241;
wire net_14121;
wire net_9106;
wire net_13653;
wire net_4070;
wire net_18256;
wire net_9327;
wire net_11173;
wire net_6272;
wire net_3141;
wire net_1670;
wire net_15939;
wire net_4274;
wire net_3265;
wire net_2801;
wire net_2932;
wire net_4951;
wire net_13342;
wire net_12420;
wire net_7928;
wire net_8277;
wire net_5812;
wire net_1264;
wire net_8077;
wire net_9852;
wire net_9300;
wire net_3148;
wire net_1229;
wire net_6316;
wire net_16148;
wire net_12746;
wire net_14385;
wire net_6277;
wire net_16125;
wire net_766;
wire net_1153;
wire net_3014;
wire net_8469;
wire net_10961;
wire net_9102;
wire net_9252;
wire net_6734;
wire net_5692;
wire net_14241;
wire x856;
wire net_18762;
wire net_18295;
wire net_3454;
wire net_5113;
wire net_9533;
wire net_13682;
wire net_12333;
wire net_3729;
wire net_10465;
wire net_18942;
wire net_14347;
wire net_9589;
wire net_2251;
wire net_12914;
wire net_8898;
wire net_9623;
wire net_7439;
wire net_10418;
wire net_9727;
wire net_955;
wire net_2585;
wire net_15670;
wire net_15952;
wire net_1996;
wire net_7046;
wire x1745;
wire net_13635;
wire net_1029;
wire net_15702;
wire net_13664;
wire net_9812;
wire net_9066;
wire net_12566;
wire net_12762;
wire net_2986;
wire net_3162;
wire net_4034;
wire net_4791;
wire net_13082;
wire net_11937;
wire net_3510;
wire net_16624;
wire net_11848;
wire net_10492;
wire net_3180;
wire net_3249;
wire net_15277;
wire net_14002;
wire net_6157;
wire net_16006;
wire net_734;
wire net_14152;
wire net_12564;
wire net_2544;
wire net_15801;
wire net_15957;
wire net_3186;
wire net_11314;
wire net_8177;
wire net_13895;
wire net_16942;
wire net_5277;
wire net_17770;
wire net_14730;
wire net_7269;
wire net_4372;
wire net_15398;
wire net_1076;
wire net_14051;
wire net_10168;
wire net_8234;
wire net_10399;
wire net_9711;
wire net_4352;
wire net_15647;
wire net_681;
wire net_7346;
wire net_18864;
wire net_13136;
wire net_6533;
wire net_5252;
wire net_17260;
wire net_146;
wire net_9562;
wire net_16250;
wire net_5752;
wire net_4594;
wire net_15009;
wire net_4454;
wire net_6290;
wire net_4624;
wire net_11522;
wire net_7621;
wire net_428;
wire net_16689;
wire net_9675;
wire net_10557;
wire net_14816;
wire net_7780;
wire net_4666;
wire net_16656;
wire net_2888;
wire net_17082;
wire net_12884;
wire net_14362;
wire net_888;
wire net_13066;
wire net_10772;
wire net_13212;
wire net_11298;
wire net_11095;
wire net_9526;
wire net_5191;
wire net_18833;
wire net_8480;
wire net_18378;
wire net_10513;
wire net_1023;
wire net_4814;
wire net_5233;
wire net_7499;
wire net_3623;
wire net_301;
wire net_2360;
wire net_3617;
wire net_7432;
wire net_1343;
wire net_18729;
wire net_7147;
wire net_2285;
wire net_16704;
wire net_12690;
wire net_7355;
wire net_16175;
wire net_16555;
wire net_590;
wire net_3879;
wire net_3240;
wire net_15150;
wire net_8229;
wire net_9342;
wire net_12135;
wire net_10094;
wire net_4194;
wire net_12361;
wire net_5464;
wire net_16136;
wire net_8335;
wire net_8530;
wire net_15059;
wire net_10145;
wire net_1736;
wire net_12807;
wire net_12258;
wire net_9814;
wire net_11660;
wire net_6947;
wire net_16363;
wire net_10314;
wire net_10574;
wire net_4148;
wire net_18854;
wire net_9155;
wire x4227;
wire net_5048;
wire net_7869;
wire net_1669;
wire net_11505;
wire net_12408;
wire net_14096;
wire net_1041;
wire net_7628;
wire net_6385;
wire net_16804;
wire net_14027;
wire net_2950;
wire net_6056;
wire net_6108;
wire net_5851;
wire net_14350;
wire net_18340;
wire net_17051;
wire net_4778;
wire net_11211;
wire net_17207;
wire net_13159;
wire net_16638;
wire net_2364;
wire net_942;
wire net_12822;
wire net_8763;
wire net_17241;
wire net_17341;
wire net_17750;
wire net_13658;
wire net_10917;
wire net_6436;
wire net_15201;
wire net_1494;
wire net_18731;
wire net_4415;
wire net_18129;
wire net_2154;
wire net_1726;
wire net_5527;
wire net_4123;
wire net_7082;
wire net_5705;
wire net_16949;
wire net_12165;
wire net_3298;
wire net_3099;
wire net_17647;
wire net_10658;
wire net_16232;
wire net_15065;
wire net_6339;
wire net_7380;
wire net_1794;
wire net_18085;
wire net_9363;
wire net_12508;
wire net_6503;
wire net_5536;
wire net_1022;
wire net_4638;
wire net_11129;
wire net_6110;
wire net_16426;
wire net_8182;
wire net_15894;
wire net_16199;
wire net_17030;
wire net_13960;
wire net_9270;
wire net_17446;
wire net_15401;
wire net_18122;
wire net_16089;
wire net_13152;
wire net_12439;
wire net_14673;
wire net_1122;
wire net_4911;
wire net_15679;
wire net_6228;
wire net_5505;
wire net_8540;
wire net_4534;
wire net_6252;
wire net_17206;
wire net_18692;
wire net_17303;
wire net_6491;
wire net_13898;
wire net_4713;
wire net_9709;
wire net_18091;
wire net_9002;
wire net_17284;
wire net_17434;
wire net_4307;
wire net_8292;
wire net_5513;
wire net_8248;
wire net_3962;
wire net_11834;
wire net_4553;
wire net_275;
wire x785;
wire net_12641;
wire net_9486;
wire net_4831;
wire net_2914;
wire net_15050;
wire net_11366;
wire net_2590;
wire net_10841;
wire net_7280;
wire net_13293;
wire net_13351;
wire net_1137;
wire net_7424;
wire net_4830;
wire net_5036;
wire net_12860;
wire net_13909;
wire net_4865;
wire net_16266;
wire net_11765;
wire net_9955;
wire net_14370;
wire net_11978;
wire net_11193;
wire net_12581;
wire net_11895;
wire net_5622;
wire net_18805;
wire net_3357;
wire net_9467;
wire net_14054;
wire net_9694;
wire net_8425;
wire net_17620;
wire net_8298;
wire net_16800;
wire x971;
wire net_14199;
wire net_14672;
wire net_943;
wire net_10413;
wire net_16736;
wire net_4392;
wire net_11330;
wire net_9435;
wire net_13088;
wire net_2542;
wire net_7594;
wire net_11996;
wire net_12537;
wire net_18035;
wire net_17009;
wire net_17642;
wire x3372;
wire net_2256;
wire net_4934;
wire net_17779;
wire net_12809;
wire net_4122;
wire net_4315;
wire net_17418;
wire net_18365;
wire net_8503;
wire net_4996;
wire net_11190;
wire net_16442;
wire net_1064;
wire net_14016;
wire net_10165;
wire net_6227;
wire net_7173;
wire net_17819;
wire net_12907;
wire net_15734;
wire net_9784;
wire net_12704;
wire net_13544;
wire net_7191;
wire net_10988;
wire net_17175;
wire net_6037;
wire net_10554;
wire net_7283;
wire net_14609;
wire net_5627;
wire net_3817;
wire net_9441;
wire net_3281;
wire net_10659;
wire net_3949;
wire net_8185;
wire net_10215;
wire net_16171;
wire net_6231;
wire net_3434;
wire net_3818;
wire net_18067;
wire net_3756;
wire net_9464;
wire net_18341;
wire net_4169;
wire net_17059;
wire net_7845;
wire net_13451;
wire net_9957;
wire net_742;
wire net_11979;
wire net_5139;
wire net_18906;
wire net_6384;
wire net_18850;
wire net_12976;
wire net_16265;
wire net_7092;
wire net_2830;
wire net_18084;
wire net_4509;
wire net_883;
wire net_11605;
wire net_13476;
wire net_8124;
wire net_4108;
wire net_2957;
wire net_9970;
wire net_446;
wire net_1712;
wire net_3063;
wire net_1499;
wire net_3295;
wire net_8242;
wire net_15060;
wire net_4379;
wire net_14985;
wire net_18943;
wire net_10000;
wire net_15141;
wire net_6114;
wire net_2303;
wire net_1735;
wire net_2210;
wire net_2176;
wire net_8249;
wire net_13191;
wire net_16592;
wire net_8563;
wire net_11933;
wire net_16130;
wire net_997;
wire net_17466;
wire net_10837;
wire net_12243;
wire net_11060;
wire net_256;
wire net_8762;
wire net_7490;
wire net_5797;
wire net_10931;
wire net_16104;
wire net_12891;
wire x4204;
wire net_4835;
wire net_16662;
wire net_5342;
wire net_7463;
wire net_11124;
wire net_13216;
wire x13786;
wire net_3987;
wire net_6557;
wire net_8468;
wire net_2219;
wire net_18418;
wire net_7343;
wire net_11166;
wire net_17264;
wire net_5680;
wire net_15657;
wire net_16176;
wire net_1876;
wire net_7483;
wire net_13130;
wire net_15567;
wire net_14611;
wire net_9810;
wire net_5116;
wire net_15218;
wire net_369;
wire net_12051;
wire net_12709;
wire net_15756;
wire net_4358;
wire net_7543;
wire net_9835;
wire net_10495;
wire net_7959;
wire net_3935;
wire net_11290;
wire net_15551;
wire net_2809;
wire net_15273;
wire net_780;
wire net_3586;
wire net_3184;
wire net_6812;
wire net_12226;
wire x12969;
wire net_15979;
wire net_9272;
wire net_10095;
wire net_5263;
wire net_155;
wire net_11350;
wire net_9301;
wire net_11357;
wire net_12555;
wire net_16553;
wire net_10636;
wire x4805;
wire net_3850;
wire net_9023;
wire net_9153;
wire net_349;
wire net_8222;
wire net_12923;
wire net_1409;
wire net_8547;
wire net_14367;
wire net_12576;
wire net_2977;
wire net_13140;
wire net_1428;
wire net_13679;
wire net_14629;
wire net_14518;
wire net_15297;
wire net_13137;
wire net_5222;
wire net_10510;
wire net_14340;
wire net_4238;
wire net_5844;
wire net_2350;
wire net_6293;
wire net_10506;
wire net_5740;
wire net_14763;
wire net_16697;
wire net_8950;
wire net_12366;
wire net_18226;
wire net_3143;
wire net_3226;
wire net_9819;
wire net_2757;
wire net_9531;
wire net_12776;
wire net_3629;
wire net_7315;
wire net_2038;
wire net_2369;
wire net_17731;
wire net_17491;
wire net_12878;
wire net_1676;
wire net_698;
wire net_14230;
wire net_12969;
wire net_14374;
wire net_5259;
wire net_17618;
wire net_8515;
wire net_4649;
wire net_2485;
wire net_6967;
wire net_13906;
wire net_3857;
wire net_18840;
wire net_749;
wire net_11729;
wire net_15053;
wire net_1948;
wire net_11500;
wire net_11898;
wire net_1006;
wire net_15922;
wire net_2781;
wire net_6767;
wire net_18264;
wire net_9724;
wire x4796;
wire net_14695;
wire net_17694;
wire net_7839;
wire net_15950;
wire net_18536;
wire net_15253;
wire net_7544;
wire net_18392;
wire net_17395;
wire net_15955;
wire net_3056;
wire net_14050;
wire net_8710;
wire net_3614;
wire net_7624;
wire net_13007;
wire net_17399;
wire net_6792;
wire net_15600;
wire net_14991;
wire net_4496;
wire net_9525;
wire net_18748;
wire net_6067;
wire net_2127;
wire net_3407;
wire net_8720;
wire net_13569;
wire net_17431;
wire net_737;
wire net_3656;
wire net_2284;
wire net_5865;
wire net_13372;
wire net_17921;
wire net_15623;
wire net_5957;
wire net_11541;
wire net_11722;
wire net_5201;
wire net_12375;
wire net_1156;
wire net_15127;
wire net_14127;
wire net_16963;
wire net_1966;
wire net_13641;
wire net_13049;
wire net_14299;
wire net_12188;
wire net_4571;
wire net_11718;
wire net_12873;
wire net_16081;
wire net_5977;
wire net_16520;
wire net_326;
wire net_2381;
wire net_10286;
wire net_11012;
wire net_17142;
wire net_15393;
wire net_9504;
wire net_5403;
wire net_15932;
wire net_10242;
wire net_6668;
wire net_6735;
wire net_3175;
wire net_10076;
wire net_14918;
wire net_17865;
wire net_2829;
wire net_10288;
wire net_3142;
wire net_4099;
wire net_4815;
wire net_1219;
wire net_12826;
wire net_14410;
wire net_10886;
wire net_10871;
wire net_13815;
wire net_3884;
wire net_2877;
wire net_3736;
wire net_8745;
wire net_9352;
wire net_8334;
wire net_1632;
wire net_3796;
wire net_1661;
wire net_1236;
wire net_13627;
wire net_8987;
wire net_13771;
wire net_19022;
wire net_2700;
wire net_18444;
wire net_17778;
wire net_7996;
wire net_7868;
wire net_10307;
wire net_16514;
wire net_9548;
wire net_17701;
wire net_1488;
wire net_6273;
wire net_6841;
wire net_2812;
wire net_15406;
wire net_352;
wire net_5691;
wire net_12721;
wire net_18140;
wire net_9320;
wire net_3920;
wire x13263;
wire net_6342;
wire net_7373;
wire net_15810;
wire net_7903;
wire net_1641;
wire net_7511;
wire x13271;
wire net_16645;
wire net_4919;
wire net_1103;
wire net_18608;
wire net_17002;
wire net_767;
wire net_16742;
wire net_4557;
wire net_9754;
wire net_5488;
wire net_8693;
wire net_2016;
wire net_4292;
wire net_7564;
wire net_14169;
wire net_17036;
wire net_7702;
wire net_10486;
wire net_16369;
wire net_3125;
wire net_13952;
wire net_10962;
wire net_12544;
wire net_6550;
wire net_18434;
wire net_9101;
wire net_13021;
wire net_9022;
wire net_19023;
wire net_10043;
wire net_15873;
wire net_16755;
wire net_13321;
wire net_7526;
wire net_14815;
wire net_468;
wire net_9308;
wire net_18916;
wire net_16433;
wire net_9257;
wire net_9372;
wire net_16596;
wire net_9738;
wire net_11654;
wire net_18077;
wire net_15573;
wire net_179;
wire net_16877;
wire net_9665;
wire net_10171;
wire net_8677;
wire net_15898;
wire net_14871;
wire net_14722;
wire net_3261;
wire net_17100;
wire net_2289;
wire net_18145;
wire net_7300;
wire net_6759;
wire net_11244;
wire net_5919;
wire net_1868;
wire net_13942;
wire net_18345;
wire net_7205;
wire net_10110;
wire net_17900;
wire net_12684;
wire net_3863;
wire net_10538;
wire net_9856;
wire net_17280;
wire net_5778;
wire net_3382;
wire net_4257;
wire net_13756;
wire net_17944;
wire net_4872;
wire net_990;
wire x3861;
wire net_7423;
wire net_11485;
wire net_11728;
wire net_10428;
wire net_10473;
wire net_11763;
wire net_3774;
wire net_1803;
wire net_13803;
wire net_8031;
wire net_1134;
wire net_363;
wire net_17025;
wire x13663;
wire net_776;
wire net_4550;
wire net_2508;
wire net_15358;
wire net_9624;
wire net_12118;
wire net_1650;
wire net_8451;
wire net_10353;
wire net_17018;
wire net_3149;
wire net_10717;
wire net_12696;
wire net_13574;
wire net_15174;
wire net_1675;
wire net_6454;
wire net_11253;
wire net_19019;
wire net_2247;
wire net_8115;
wire net_2291;
wire net_6525;
wire net_10531;
wire net_11108;
wire net_15220;
wire net_16045;
wire net_11096;
wire net_15558;
wire net_8414;
wire net_18802;
wire net_1201;
wire net_2525;
wire net_12404;
wire net_12073;
wire net_9701;
wire net_14331;
wire net_5106;
wire net_8074;
wire net_13852;
wire net_859;
wire net_1167;
wire net_7259;
wire net_8636;
wire net_1044;
wire net_18561;
wire net_4322;
wire net_10948;
wire net_10617;
wire net_2043;
wire net_18609;
wire net_6775;
wire net_10662;
wire net_15818;
wire net_3605;
wire net_14336;
wire net_6635;
wire net_10865;
wire net_12174;
wire net_4114;
wire net_7250;
wire net_11055;
wire net_17425;
wire net_14220;
wire net_865;
wire net_10330;
wire net_13500;
wire net_9896;
wire net_2621;
wire net_13326;
wire net_13832;
wire net_1223;
wire net_2750;
wire net_5816;
wire net_926;
wire net_11961;
wire net_4623;
wire net_7264;
wire x4693;
wire net_7403;
wire net_17654;
wire net_6153;
wire net_14656;
wire net_8642;
wire net_7188;
wire net_10595;
wire net_12868;
wire net_9185;
wire net_6466;
wire net_2048;
wire net_18471;
wire net_4481;
wire net_3633;
wire net_7337;
wire net_7036;
wire net_14705;
wire net_3561;
wire net_1295;
wire net_1543;
wire net_10993;
wire net_13692;
wire net_9429;
wire net_5661;
wire net_2071;
wire net_1923;
wire net_1275;
wire net_13481;
wire net_11031;
wire net_13463;
wire net_940;
wire net_4411;
wire net_3719;
wire net_4857;
wire net_10572;
wire net_15681;
wire net_6061;
wire net_8311;
wire net_5350;
wire net_12330;
wire net_14329;
wire net_9627;
wire net_13631;
wire net_5335;
wire net_12849;
wire net_18578;
wire net_19035;
wire net_10133;
wire net_12438;
wire net_9485;
wire net_16786;
wire net_17503;
wire net_1454;
wire net_6949;
wire net_17793;
wire net_3342;
wire net_14711;
wire net_1550;
wire net_9642;
wire net_10069;
wire net_233;
wire net_18596;
wire net_5138;
wire net_18629;
wire net_3459;
wire net_16154;
wire net_13411;
wire net_1268;
wire net_11127;
wire net_3780;
wire net_13783;
wire net_1115;
wire net_4051;
wire net_11465;
wire net_17820;
wire net_6641;
wire net_961;
wire net_18886;
wire net_9643;
wire net_2106;
wire net_14691;
wire net_5175;
wire net_11909;
wire net_14196;
wire net_4894;
wire x13654;
wire net_9424;
wire net_3327;
wire net_9480;
wire net_5091;
wire net_18189;
wire net_13719;
wire net_3456;
wire net_13700;
wire net_7627;
wire net_12250;
wire net_12453;
wire net_13220;
wire net_9907;
wire net_4407;
wire net_13713;
wire net_16485;
wire net_1586;
wire net_14113;
wire net_5354;
wire net_216;
wire net_13284;
wire net_10727;
wire net_18667;
wire net_2881;
wire net_12630;
wire net_4602;
wire x105;
wire net_15556;
wire net_12057;
wire net_5635;
wire net_9495;
wire net_16198;
wire net_8379;
wire net_8806;
wire net_11237;
wire net_9097;
wire net_12520;
wire net_1120;
wire net_5881;
wire net_2848;
wire net_7126;
wire net_973;
wire net_11832;
wire net_1139;
wire net_6998;
wire net_7394;
wire net_9337;
wire net_3902;
wire net_18291;
wire net_1574;
wire x1305;
wire net_9008;
wire net_4842;
wire net_11576;
wire net_154;
wire net_8016;
wire net_3699;
wire net_16796;
wire net_13847;
wire net_12056;
wire net_14946;
wire net_1478;
wire net_14075;
wire net_587;
wire net_1696;
wire net_2179;
wire net_1262;
wire net_9163;
wire net_17892;
wire net_4027;
wire net_14106;
wire net_8750;
wire net_4213;
wire net_4505;
wire net_18170;
wire net_17517;
wire net_4131;
wire net_7396;
wire net_10779;
wire net_14937;
wire net_1907;
wire net_11323;
wire net_18898;
wire net_16201;
wire net_15420;
wire net_16982;
wire net_4164;
wire net_6312;
wire net_195;
wire net_10200;
wire net_18663;
wire net_10247;
wire net_16110;
wire net_10104;
wire net_17093;
wire net_8980;
wire net_13999;
wire net_18891;
wire net_8323;
wire net_9042;
wire net_7002;
wire net_3761;
wire net_9196;
wire net_13722;
wire net_242;
wire net_7076;
wire net_7719;
wire net_7722;
wire x4932;
wire net_18724;
wire net_9543;
wire net_8938;
wire net_11384;
wire net_8336;
wire net_13514;
wire net_1311;
wire net_5939;
wire net_11230;
wire net_13307;
wire net_7068;
wire net_10207;
wire net_18732;
wire net_10549;
wire net_11911;
wire net_17278;
wire x13440;
wire net_5937;
wire net_8208;
wire net_12314;
wire net_3558;
wire net_9678;
wire net_555;
wire net_16327;
wire net_1613;
wire net_7758;
wire net_13016;
wire net_15051;
wire net_790;
wire net_11938;
wire net_14665;
wire net_1417;
wire net_11466;
wire net_18501;
wire net_11520;
wire net_13423;
wire net_2386;
wire net_11063;
wire net_2166;
wire net_8359;
wire net_11588;
wire net_17918;
wire net_12830;
wire net_15846;
wire net_10650;
wire net_7150;
wire net_13699;
wire net_6537;
wire net_14873;
wire net_17497;
wire net_4416;
wire net_714;
wire net_5015;
wire net_1309;
wire net_2999;
wire net_9567;
wire net_683;
wire net_1771;
wire net_148;
wire net_4493;
wire net_12136;
wire net_13555;
wire net_7220;
wire net_17544;
wire net_9171;
wire net_17950;
wire net_15852;
wire net_7449;
wire net_7751;
wire net_10362;
wire net_15799;
wire net_14504;
wire net_5547;
wire net_9361;
wire net_15411;
wire net_9149;
wire net_5616;
wire net_7353;
wire net_12117;
wire net_7113;
wire net_8588;
wire net_2403;
wire net_7740;
wire net_15173;
wire net_17957;
wire net_15582;
wire net_14147;
wire net_7913;
wire net_15238;
wire net_18828;
wire net_16220;
wire net_8550;
wire net_14761;
wire net_16819;
wire net_394;
wire net_810;
wire net_1548;
wire net_15861;
wire net_17159;
wire net_1189;
wire net_3778;
wire net_409;
wire net_7183;
wire net_15366;
wire net_3470;
wire net_11908;
wire net_16297;
wire net_13354;
wire net_8036;
wire net_16790;
wire net_18393;
wire net_11509;
wire net_15113;
wire net_3419;
wire net_10754;
wire net_16021;
wire net_17807;
wire net_1254;
wire net_10733;
wire net_11417;
wire net_18708;
wire net_15616;
wire net_12793;
wire net_13171;
wire net_10533;
wire net_7240;
wire net_11862;
wire net_7365;
wire net_5361;
wire x912;
wire net_15496;
wire net_8703;
wire net_9383;
wire net_9841;
wire net_4675;
wire net_8378;
wire net_327;
wire net_3877;
wire net_16139;
wire net_16583;
wire net_353;
wire net_8052;
wire net_13799;
wire net_11730;
wire net_12322;
wire net_9584;
wire x764;
wire net_8552;
wire net_16620;
wire net_5730;
wire net_14209;
wire net_8770;
wire net_14140;
wire net_6927;
wire net_12628;
wire net_3046;
wire net_164;
wire net_6019;
wire net_4702;
wire net_7632;
wire net_15396;
wire net_17583;
wire net_3096;
wire net_1629;
wire net_8947;
wire net_14950;
wire net_11387;
wire net_14431;
wire net_805;
wire net_3277;
wire net_12032;
wire net_6740;
wire net_12093;
wire net_3590;
wire net_2151;
wire net_17198;
wire net_8521;
wire net_2688;
wire net_14304;
wire net_1622;
wire net_13392;
wire net_5149;
wire net_6299;
wire net_11664;
wire net_16003;
wire net_17635;
wire net_7815;
wire x13291;
wire net_7453;
wire net_14793;
wire net_12998;
wire net_11744;
wire net_13420;
wire net_18685;
wire net_2244;
wire net_12825;
wire net_15809;
wire net_11737;
wire net_7826;
wire net_783;
wire net_11955;
wire net_13686;
wire net_9211;
wire net_6305;
wire net_11703;
wire net_17549;
wire net_2605;
wire net_9469;
wire net_550;
wire net_9875;
wire net_10821;
wire net_5238;
wire net_12292;
wire net_17759;
wire net_9158;
wire net_3991;
wire net_5086;
wire net_10912;
wire net_461;
wire net_14516;
wire net_7778;
wire net_16517;
wire net_6879;
wire net_12962;
wire net_6657;
wire net_8524;
wire net_9284;
wire net_14185;
wire net_1512;
wire net_17744;
wire net_18636;
wire net_15370;
wire net_14593;
wire net_8047;
wire net_1330;
wire net_5025;
wire net_4275;
wire net_17586;
wire net_3015;
wire net_11011;
wire net_1785;
wire net_4771;
wire net_11077;
wire net_13507;
wire net_16062;
wire net_17132;
wire net_10680;
wire net_9516;
wire net_6870;
wire net_16752;
wire net_9655;
wire net_5060;
wire x394;
wire net_12596;
wire net_15848;
wire net_5668;
wire net_10408;
wire net_985;
wire net_4679;
wire net_16492;
wire net_6719;
wire net_12190;
wire net_7061;
wire net_15494;
wire net_16609;
wire net_424;
wire net_6837;
wire net_1729;
wire net_3353;
wire net_12623;
wire net_16274;
wire net_4247;
wire net_17477;
wire net_5719;
wire net_17112;
wire net_3639;
wire net_14404;
wire net_15915;
wire net_8065;
wire net_12311;
wire net_12148;
wire net_11992;
wire net_3086;
wire net_4585;
wire net_2058;
wire net_11110;
wire net_3045;
wire net_12206;
wire net_17669;
wire net_4875;
wire net_2018;
wire net_13100;
wire net_11731;
wire net_2510;
wire net_9952;
wire net_3808;
wire net_7881;
wire net_12941;
wire net_14631;
wire net_6243;
wire net_7882;
wire net_6415;
wire net_14393;
wire net_18316;
wire net_9201;
wire net_17666;
wire net_6302;
wire net_8916;
wire net_2279;
wire net_14048;
wire net_3447;
wire net_15633;
wire net_6174;
wire net_8401;
wire net_14588;
wire net_17812;
wire x845;
wire x13047;
wire net_18487;
wire net_17408;
wire net_17224;
wire net_9267;
wire net_10826;
wire net_13893;
wire net_8497;
wire net_18284;
wire net_17521;
wire net_10295;
wire net_7801;
wire net_3217;
wire net_1291;
wire net_4387;
wire net_6362;
wire net_1865;
wire net_13896;
wire net_18695;
wire net_5168;
wire net_6076;
wire x2494;
wire net_5329;
wire net_18312;
wire net_14541;
wire net_10985;
wire net_17752;
wire net_8460;
wire net_10490;
wire net_2578;
wire net_8658;
wire net_16392;
wire net_1433;
wire net_10462;
wire net_18052;
wire net_17042;
wire net_11672;
wire net_13745;
wire net_15503;
wire net_14786;
wire net_8606;
wire net_5440;
wire net_9425;
wire net_2574;
wire net_5928;
wire x12962;
wire net_14235;
wire net_3531;
wire net_3747;
wire x649;
wire net_18454;
wire net_5732;
wire net_12212;
wire net_8593;
wire net_18594;
wire net_1844;
wire net_389;
wire net_11512;
wire net_902;
wire net_13981;
wire net_11287;
wire net_15859;
wire net_15907;
wire net_13237;
wire net_736;
wire net_8771;
wire net_5462;
wire net_5282;
wire net_6498;
wire net_8372;
wire net_18767;
wire net_15737;
wire net_6262;
wire net_17713;
wire net_10905;
wire net_15379;
wire net_19005;
wire net_12517;
wire net_18400;
wire x3079;
wire net_14092;
wire net_10034;
wire net_7249;
wire net_18137;
wire net_15152;
wire net_5717;
wire net_869;
wire net_3714;
wire net_12144;
wire net_8308;
wire net_11280;
wire net_4077;
wire net_2441;
wire net_18825;
wire net_4749;
wire net_5828;
wire net_6799;
wire net_8775;
wire net_12092;
wire net_13774;
wire net_2459;
wire net_15512;
wire net_10394;
wire net_14434;
wire net_5422;
wire net_6629;
wire net_6704;
wire net_12395;
wire net_15329;
wire net_19002;
wire x4420;
wire net_16415;
wire net_6508;
wire net_15832;
wire net_18968;
wire net_2075;
wire net_2548;
wire net_3359;
wire net_5848;
wire net_15883;
wire net_10085;
wire net_12296;
wire net_9069;
wire net_15900;
wire net_7548;
wire net_12889;
wire net_14866;
wire net_6165;
wire net_4795;
wire net_511;
wire net_9263;
wire net_12759;
wire net_3967;
wire net_2654;
wire net_1819;
wire net_2911;
wire net_11791;
wire net_8258;
wire net_15509;
wire net_12821;
wire net_12763;
wire net_17404;
wire net_7236;
wire net_17271;
wire net_11379;
wire net_13181;
wire net_9031;
wire net_18508;
wire net_13661;
wire net_11083;
wire net_989;
wire net_8446;
wire net_17629;
wire net_458;
wire net_18512;
wire net_11748;
wire net_7442;
wire net_8322;
wire net_14471;
wire net_9030;
wire net_10998;
wire net_16686;
wire net_10957;
wire net_14183;
wire net_13333;
wire net_4616;
wire net_11408;
wire net_13096;
wire net_16186;
wire net_4786;
wire net_16212;
wire net_8616;
wire net_18779;
wire net_5893;
wire net_7872;
wire net_10542;
wire net_17287;
wire net_10891;
wire net_2111;
wire net_3410;
wire net_14954;
wire net_5525;
wire net_8162;
wire net_12496;
wire net_16867;
wire x3874;
wire x4919;
wire net_5610;
wire net_14894;
wire x13742;
wire net_16627;
wire net_14278;
wire net_13045;
wire net_2535;
wire net_3191;
wire net_13165;
wire net_13822;
wire net_14396;
wire net_15106;
wire net_10355;
wire net_12865;
wire net_18093;
wire net_12125;
wire net_2983;
wire net_12916;
wire net_14617;
wire net_10024;
wire net_1647;
wire net_198;
wire net_12460;
wire net_10058;
wire net_7509;
wire net_4756;
wire net_5196;
wire net_13280;
wire net_15293;
wire net_16255;
wire x4036;
wire net_18476;
wire net_2892;
wire net_13263;
wire net_15646;
wire net_18711;
wire net_13077;
wire net_4444;
wire net_848;
wire net_9550;
wire net_1080;
wire net_12022;
wire net_10641;
wire net_16705;
wire net_1890;
wire net_13648;
wire net_18755;
wire net_11293;
wire net_2357;
wire net_4501;
wire net_12449;
wire net_13319;
wire net_11114;
wire net_18736;
wire net_5492;
wire net_11772;
wire net_17875;
wire net_12383;
wire net_11372;
wire net_10199;
wire net_6536;
wire net_15728;
wire net_4363;
wire net_7417;
wire net_606;
wire net_16016;
wire net_623;
wire net_3906;
wire net_663;
wire net_12503;
wire net_1891;
wire net_5180;
wire net_579;
wire net_3998;
wire net_16443;
wire net_9490;
wire net_8597;
wire net_2062;
wire net_18074;
wire net_13666;
wire net_9828;
wire net_18380;
wire net_6418;
wire net_10844;
wire net_17678;
wire net_4834;
wire net_7296;
wire net_17673;
wire net_8061;
wire net_9317;
wire net_4067;
wire net_4717;
wire net_1518;
wire net_17682;
wire net_4618;
wire net_1437;
wire net_1194;
wire net_18273;
wire net_15837;
wire net_5517;
wire net_17576;
wire net_17150;
wire net_6770;
wire net_7587;
wire net_11923;
wire net_1664;
wire net_17345;
wire net_13651;
wire net_15718;
wire net_16227;
wire net_705;
wire net_10326;
wire net_2948;
wire net_10523;
wire net_17055;
wire net_1036;
wire net_18186;
wire net_5608;
wire net_6052;
wire net_7497;
wire net_11966;
wire net_4537;
wire net_1196;
wire net_3973;
wire net_6331;
wire x2542;
wire net_6762;
wire net_9077;
wire net_5531;
wire net_6085;
wire net_6598;
wire net_5701;
wire net_11786;
wire net_3136;
wire net_4090;
wire net_12553;
wire net_6149;
wire net_9178;
wire net_10809;
wire net_3834;
wire net_10300;
wire net_13471;
wire net_3152;
wire net_14311;
wire net_3648;
wire net_1722;
wire net_16854;
wire net_2008;
wire net_6395;
wire net_18133;
wire net_11633;
wire net_2808;
wire net_18481;
wire net_8265;
wire net_9055;
wire net_14008;
wire net_17761;
wire net_6575;
wire net_16907;
wire net_16654;
wire net_4707;
wire net_6432;
wire net_13918;
wire net_16119;
wire net_17932;
wire net_957;
wire net_12771;
wire net_15667;
wire net_18839;
wire net_1287;
wire net_10625;
wire net_14040;
wire net_2726;
wire net_1340;
wire net_7277;
wire net_7165;
wire net_9599;
wire x2948;
wire net_12363;
wire net_2844;
wire net_12415;
wire net_9977;
wire net_5538;
wire net_4852;
wire net_6804;
wire net_9941;
wire net_10341;
wire net_14361;
wire net_4437;
wire net_10435;
wire net_18281;
wire net_4028;
wire net_2860;
wire net_432;
wire net_4927;
wire net_6025;
wire net_6329;
wire net_10627;
wire net_1142;
wire net_14556;
wire net_3159;
wire x13086;
wire net_5644;
wire net_16380;
wire net_2240;
wire net_14600;
wire net_18859;
wire net_2416;
wire net_12882;
wire net_6404;
wire net_8727;
wire net_14354;
wire net_6185;
wire net_9713;
wire net_5383;
wire net_17833;
wire net_10540;
wire net_7487;
wire net_13520;
wire net_4013;
wire net_11517;
wire net_2144;
wire net_2236;
wire net_11057;
wire net_3443;
wire net_3945;
wire net_8824;
wire x852;
wire net_11529;
wire net_14622;
wire net_1505;
wire net_16476;
wire net_8279;
wire net_13836;
wire net_3669;
wire net_3952;
wire net_1861;
wire net_13448;
wire net_9999;
wire net_4388;
wire net_11852;
wire net_1594;
wire net_221;
wire net_5672;
wire net_18252;
wire net_542;
wire net_14218;
wire net_17872;
wire net_13026;
wire net_12483;
wire net_6487;
wire net_18818;
wire x13494;
wire net_4562;
wire net_9437;
wire net_2376;
wire net_1520;
wire net_6562;
wire net_6713;
wire net_18529;
wire net_15867;
wire net_16767;
wire net_8579;
wire net_9638;
wire net_16619;
wire net_15287;
wire net_8005;
wire net_3664;
wire net_3233;
wire net_5124;
wire net_14521;
wire net_9731;
wire net_16642;
wire net_7178;
wire net_10937;
wire net_17212;
wire net_11814;
wire net_9649;
wire net_1584;
wire net_16693;
wire net_13539;
wire net_12612;
wire net_2330;
wire net_7890;
wire net_3397;
wire net_16348;
wire net_9777;
wire net_5898;
wire net_18976;
wire net_6785;
wire net_15948;
wire net_4391;
wire net_7814;
wire net_11473;
wire net_9045;
wire net_12659;
wire net_6875;
wire net_2857;
wire net_8674;
wire net_2767;
wire net_9594;
wire net_6120;
wire net_16837;
wire net_11491;
wire net_6604;
wire net_12652;
wire net_825;
wire net_309;
wire net_18522;
wire net_1366;
wire net_17185;
wire net_13054;
wire net_2615;
wire net_14978;
wire net_14268;
wire net_9290;
wire net_16313;
wire net_7367;
wire net_8158;
wire net_1151;
wire net_16120;
wire x838;
wire net_5240;
wire net_5318;
wire net_9993;
wire net_11138;
wire net_17149;
wire net_8291;
wire net_15046;
wire net_2818;
wire net_3213;
wire net_7690;
wire net_580;
wire net_4173;
wire net_2136;
wire net_9805;
wire net_2339;
wire net_7699;
wire net_8884;
wire net_4157;
wire net_1879;
wire net_14821;
wire net_6663;
wire net_12122;
wire net_13224;
wire net_8202;
wire net_4221;
wire net_4941;
wire net_17447;
wire net_6732;
wire net_12524;
wire net_12683;
wire net_17047;
wire net_5604;
wire net_11022;
wire net_11612;
wire net_8351;
wire net_18922;
wire net_4887;
wire net_15760;
wire net_18012;
wire net_13116;
wire net_763;
wire net_13704;
wire net_16285;
wire net_14088;
wire net_7762;
wire net_1740;
wire net_5639;
wire net_14495;
wire net_17217;
wire net_9455;
wire net_872;
wire net_9125;
wire net_10502;
wire net_8251;
wire net_3880;
wire net_5581;
wire net_18110;
wire net_16405;
wire net_4333;
wire net_11285;
wire net_14776;
wire net_18989;
wire net_5558;
wire net_7575;
wire net_4880;
wire net_1812;
wire net_8174;
wire net_12584;
wire net_4825;
wire net_10850;
wire net_18604;
wire net_8696;
wire net_4138;
wire net_3203;
wire net_12811;
wire net_11881;
wire net_2589;
wire net_2659;
wire net_7515;
wire net_12670;
wire net_591;
wire net_1700;
wire net_12739;
wire net_12985;
wire net_16766;
wire net_7557;
wire net_10188;
wire net_178;
wire net_18813;
wire net_18794;
wire net_11751;
wire net_15266;
wire net_9074;
wire net_2843;
wire net_6780;
wire net_14081;
wire net_7961;
wire net_10191;
wire net_15322;
wire net_3807;
wire net_10480;
wire net_809;
wire net_13995;
wire net_8393;
wire net_635;
wire net_1235;
wire net_266;
wire net_4279;
wire net_2691;
wire net_18041;
wire net_8610;
wire net_12600;
wire net_6622;
wire net_6007;
wire net_15520;
wire net_13205;
wire net_10176;
wire net_6549;
wire net_6542;
wire net_3460;
wire net_13091;
wire net_12859;
wire net_18811;
wire net_3198;
wire net_1626;
wire net_5720;
wire net_8366;
wire net_2822;
wire net_7317;
wire net_1258;
wire net_8413;
wire net_17857;
wire net_12041;
wire net_9866;
wire net_318;
wire net_10231;
wire net_3927;
wire net_10859;
wire net_1971;
wire net_8931;
wire net_2409;
wire net_1900;
wire net_3192;
wire net_1779;
wire net_2647;
wire net_5218;
wire net_8492;
wire net_7972;
wire net_228;
wire net_11886;
wire net_4737;
wire net_2640;
wire net_966;
wire net_13011;
wire net_7083;
wire net_3372;
wire net_4698;
wire net_2201;
wire net_6049;
wire net_2025;
wire net_2827;
wire net_16748;
wire net_2936;
wire net_7905;
wire net_5643;
wire net_9936;
wire net_5728;
wire net_13736;
wire net_16760;
wire net_17507;
wire net_8013;
wire net_17146;
wire net_10702;
wire net_12425;
wire net_10366;
wire net_16924;
wire net_14297;
wire net_11414;
wire net_10920;
wire net_11265;
wire net_12444;
wire net_15024;
wire net_12529;
wire net_10579;
wire net_16536;
wire net_7997;
wire x451;
wire net_4522;
wire net_11925;
wire net_8908;
wire net_14836;
wire net_3652;
wire net_8689;
wire net_2669;
wire net_6829;
wire net_18929;
wire net_4083;
wire net_1173;
wire net_1754;
wire net_2328;
wire net_7715;
wire net_11401;
wire net_16561;
wire net_8080;
wire net_5571;
wire net_15302;
wire net_5805;
wire net_10205;
wire net_12792;
wire net_7254;
wire net_13623;
wire net_7684;
wire net_17607;
wire net_16164;
wire net_12991;
wire net_10743;
wire net_9604;
wire net_13565;
wire net_13605;
wire net_14467;
wire net_6887;
wire net_18263;
wire net_9838;
wire net_15427;
wire net_4462;
wire net_15546;
wire net_11038;
wire net_1394;
wire net_2963;
wire net_5412;
wire net_5546;
wire net_6134;
wire net_1281;
wire net_9395;
wire net_2463;
wire net_9291;
wire net_8210;
wire net_15945;
wire net_16996;
wire net_8995;
wire net_11258;
wire net_8367;
wire net_4058;
wire net_8432;
wire net_16469;
wire net_3509;
wire net_1162;
wire net_13856;
wire net_17536;
wire net_2472;
wire net_2742;
wire net_2790;
wire net_13589;
wire net_13120;
wire net_5007;
wire net_10738;
wire net_10318;
wire net_15386;
wire net_10434;
wire net_13795;
wire net_8360;
wire net_11902;
wire net_6521;
wire net_10269;
wire net_17480;
wire x13605;
wire net_3320;
wire net_10561;
wire net_17599;
wire net_16108;
wire net_5221;
wire net_3657;
wire net_5550;
wire net_1353;
wire net_14683;
wire net_11652;
wire net_15165;
wire net_5303;
wire net_3581;
wire net_18932;
wire net_14961;
wire net_4049;
wire net_1300;
wire net_18876;
wire net_18644;
wire net_14322;
wire net_12131;
wire net_16723;
wire net_14419;
wire net_16102;
wire net_17312;
wire net_13432;
wire net_547;
wire net_10941;
wire net_14026;
wire net_1098;
wire net_10049;
wire net_6683;
wire net_238;
wire net_3074;
wire net_5475;
wire net_8973;
wire net_7055;
wire net_11354;
wire net_2438;
wire net_7896;
wire net_1911;
wire net_6906;
wire net_17512;
wire net_649;
wire net_13597;
wire net_1374;
wire net_13887;
wire net_4843;
wire net_8959;
wire net_16887;
wire net_2494;
wire net_18671;
wire net_15747;
wire net_11217;
wire net_16989;
wire net_6819;
wire net_12274;
wire net_14811;
wire net_3700;
wire net_13349;
wire net_530;
wire net_9140;
wire net_15155;
wire net_10529;
wire net_11839;
wire net_10004;
wire net_673;
wire net_4268;
wire net_7022;
wire net_7029;
wire net_12247;
wire net_2797;
wire net_6256;
wire net_9966;
wire net_3846;
wire net_12261;
wire net_3549;
wire net_9790;
wire net_1445;
wire net_8581;
wire net_10227;
wire net_6729;
wire net_13807;
wire net_16206;
wire net_9922;
wire net_7639;
wire net_10126;
wire net_11454;
wire net_11583;
wire net_5379;
wire net_13340;
wire net_3913;
wire x827;
wire net_9988;
wire net_11643;
wire net_3787;
wire net_17487;
wire net_1810;
wire net_1118;
wire net_10776;
wire net_372;
wire net_6858;
wire net_12235;
wire net_9882;
wire net_18678;
wire net_7086;
wire net_2990;
wire net_6324;
wire net_16145;
wire net_11749;
wire net_18741;
wire net_3595;
wire net_2788;
wire net_8923;
wire net_10383;
wire net_13787;
wire net_6899;
wire net_10142;
wire net_14490;
wire net_15774;
wire x20;
wire net_3489;
wire net_15346;
wire net_11184;
wire net_19047;
wire net_13581;
wire net_563;
wire net_7854;
wire net_1147;
wire net_13979;
wire net_18194;
wire net_13388;
wire net_15242;
wire net_15193;
wire net_8815;
wire net_13452;
wire net_2158;
wire net_4366;
wire net_10234;
wire net_10175;
wire net_13936;
wire net_17997;
wire net_5009;
wire net_12254;
wire net_3684;
wire net_14677;
wire net_8418;
wire x76;
wire net_2428;
wire net_10695;
wire net_8652;
wire net_10814;
wire net_2895;
wire net_13299;
wire net_15488;
wire net_15985;
wire net_8238;
wire net_13418;
wire net_2477;
wire net_12957;
wire net_9927;
wire net_16238;
wire net_5653;
wire net_13819;
wire net_16770;
wire net_7664;
wire net_4188;
wire net_15451;
wire net_4040;
wire net_6146;
wire net_5433;
wire net_12766;
wire net_3759;
wire net_3511;
wire net_374;
wire net_12839;
wire net_14069;
wire net_8755;
wire net_17076;
wire net_1987;
wire net_12816;
wire net_16242;
wire net_12910;
wire net_7011;
wire net_249;
wire net_3602;
wire net_16827;
wire net_13155;
wire net_17258;
wire net_9963;
wire net_17122;
wire net_5283;
wire net_18215;
wire net_9013;
wire net_8871;
wire net_15895;
wire net_6196;
wire net_4009;
wire net_10766;
wire net_13488;
wire net_17937;
wire net_7648;
wire net_8508;
wire net_13880;
wire net_5993;
wire net_2632;
wire net_16028;
wire net_2547;
wire net_5076;
wire net_8634;
wire net_16487;
wire x4448;
wire net_17167;
wire net_9084;
wire net_15440;
wire net_2295;
wire net_5831;
wire net_5628;
wire net_1817;
wire net_17962;
wire net_11009;
wire net_9348;
wire net_16078;
wire net_1381;
wire net_6445;
wire net_202;
wire net_3312;
wire net_13596;
wire net_17590;
wire net_1756;
wire net_7325;
wire net_18491;
wire net_2208;
wire net_6475;
wire net_918;
wire net_7727;
wire net_11204;
wire net_5397;
wire net_18573;
wire net_9204;
wire net_17374;
wire net_5901;
wire net_13610;
wire net_9356;
wire net_1129;
wire net_10780;
wire net_1056;
wire net_11345;
wire net_14689;
wire net_4908;
wire net_14561;
wire net_10896;
wire net_17969;
wire net_4781;
wire net_2044;
wire net_17458;
wire net_2181;
wire net_7402;
wire net_6913;
wire net_8626;
wire net_14782;
wire net_18414;
wire net_8406;
wire net_17508;
wire net_4530;
wire net_7379;
wire net_838;
wire net_6123;
wire net_10441;
wire net_18303;
wire net_16899;
wire net_11151;
wire net_14316;
wire net_14202;
wire x4192;
wire net_11750;
wire net_5872;
wire net_4980;
wire net_7107;
wire net_17846;
wire net_11270;
wire net_15341;
wire net_3827;
wire net_16542;
wire net_8405;
wire net_12072;
wire net_5308;
wire net_3515;
wire net_5033;
wire net_12747;
wire net_16059;
wire net_8085;
wire net_17171;
wire net_9720;
wire net_18153;
wire net_3398;
wire net_9223;
wire net_16721;
wire net_342;
wire net_13400;
wire net_612;
wire net_892;
wire net_16930;
wire net_8098;
wire net_4198;
wire net_12871;
wire net_10423;
wire net_5434;
wire net_11144;
wire net_10848;
wire net_14488;
wire net_8344;
wire net_12639;
wire net_6511;
wire net_10060;
wire net_1537;
wire net_11105;
wire net_13051;
wire net_13399;
wire net_4074;
wire net_16730;
wire net_4000;
wire net_2214;
wire net_14913;
wire net_3338;
wire net_16073;
wire net_17973;
wire net_5987;
wire net_15468;
wire net_13238;
wire net_417;
wire net_9929;
wire net_17370;
wire net_5387;
wire net_10634;
wire net_8217;
wire x13863;
wire net_7467;
wire net_10758;
wire net_17191;
wire net_17011;
wire net_3337;
wire net_8287;
wire net_2662;
wire net_3752;
wire net_482;
wire net_5144;
wire net_10805;
wire net_3258;
wire net_10942;
wire x552;
wire net_149;
wire net_15437;
wire net_7790;
wire net_13107;
wire net_13127;
wire x1195;
wire net_5160;
wire net_15995;
wire net_6494;
wire net_14137;
wire x13619;
wire net_15035;
wire net_577;
wire net_3401;
wire net_13245;
wire net_10313;
wire net_2550;
wire net_797;
wire net_7747;
wire net_3545;
wire net_1799;
wire net_10150;
wire net_11224;
wire net_15132;
wire net_11859;
wire net_16092;
wire net_18544;
wire net_9218;
wire net_12909;
wire net_337;
wire net_10581;
wire net_13312;
wire net_4476;
wire net_690;
wire net_17729;
wire net_6820;
wire net_7933;
wire net_3743;
wire net_523;
wire net_11070;
wire net_6718;
wire net_7144;
wire net_3375;
wire net_6744;
wire net_9620;
wire net_18620;
wire net_4926;
wire net_3467;
wire net_16637;
wire net_9617;
wire net_15785;
wire net_8972;
wire net_9760;
wire net_17243;
wire net_16439;
wire net_4467;
wire net_12129;
wire net_5028;
wire net_4721;
wire net_18179;
wire net_5756;
wire net_18999;
wire net_1631;
wire net_4426;
wire net_16955;
wire net_1337;
wire net_5786;
wire net_1182;
wire net_14254;
wire net_17768;
wire net_7231;
wire net_16286;
wire net_13656;
wire net_14458;
wire net_18244;
wire net_1950;
wire net_9052;
wire net_15067;
wire net_18973;
wire x13031;
wire net_9280;
wire net_7039;
wire net_14803;
wire net_2421;
wire net_5684;
wire net_4901;
wire net_4804;
wire net_880;
wire net_1402;
wire net_18784;
wire net_18337;
wire net_4100;
wire net_18028;
wire net_8474;
wire net_17470;
wire net_16600;
wire net_8535;
wire x13612;
wire net_5151;
wire net_16309;
wire net_13922;
wire net_2901;
wire net_11876;
wire net_15792;
wire net_4950;
wire net_13255;
wire net_4944;
wire net_18103;
wire net_18298;
wire net_4847;
wire net_12661;
wire net_3052;
wire net_6652;
wire net_10906;
wire net_7295;
wire net_11554;
wire net_6368;
wire net_16939;
wire net_14889;
wire net_487;
wire net_7992;
wire net_8861;
wire net_17785;
wire net_5056;
wire net_756;
wire net_7735;
wire net_13636;
wire net_4765;
wire net_17614;
wire net_14234;
wire net_7798;
wire net_10101;
wire net_12230;
wire net_17841;
wire net_5031;
wire net_11301;
wire net_15477;
wire net_17319;
wire net_17724;
wire net_11845;
wire net_3537;
wire net_18447;
wire net_15541;
wire net_12897;
wire net_2225;
wire net_7659;
wire net_16356;
wire net_16342;
wire net_17104;
wire net_16917;
wire net_15257;
wire net_4741;
wire net_11687;
wire net_16334;
wire net_15720;
wire net_9402;
wire net_10469;
wire net_12852;
wire net_16501;
wire net_11420;
wire x668;
wire net_174;
wire net_7987;
wire net_7214;
wire net_15208;
wire net_1831;
wire net_6202;
wire net_11691;
wire net_1482;
wire net_17600;
wire net_3291;
wire net_2928;
wire net_3306;
wire net_14573;
wire net_17829;
wire net_7563;
wire net_14460;
wire net_1485;
wire net_4129;
wire net_9236;
wire net_10272;
wire net_10053;
wire net_3245;
wire net_13300;
wire net_16902;
wire net_9385;
wire net_7473;
wire x208;
wire net_6920;
wire net_7335;
wire net_14742;
wire net_7387;
wire net_11987;
wire net_10787;
wire net_12711;
wire net_12740;
wire net_13407;
wire net_13929;
wire net_745;
wire net_9651;
wire net_14737;
wire net_17774;
wire net_16352;
wire net_14271;
wire net_1244;
wire net_15919;
wire net_429;
wire net_10966;
wire net_12593;
wire net_356;
wire net_13701;
wire net_545;
wire net_11432;
wire net_2147;
wire net_11700;
wire net_10361;
wire net_560;
wire net_9253;
wire net_10098;
wire net_5148;
wire net_4603;
wire net_15120;
wire net_14017;
wire net_17705;
wire net_15586;
wire net_17984;
wire net_5510;
wire net_11951;
wire net_9359;
wire net_10500;
wire net_6709;
wire net_7310;
wire net_16874;
wire net_13151;
wire net_7522;
wire net_2872;
wire net_2432;
wire net_6833;
wire net_12780;
wire net_5401;
wire net_322;
wire net_420;
wire net_2322;
wire net_8944;
wire net_4344;
wire net_9109;
wire x3968;
wire net_3341;
wire net_13376;
wire net_1072;
wire net_7136;
wire net_13738;
wire net_18737;
wire net_15527;
wire net_4510;
wire net_11113;
wire net_19014;
wire net_6278;
wire net_1730;
wire net_6311;
wire net_4575;
wire net_13501;
wire net_651;
wire net_15766;
wire net_18370;
wire net_14653;
wire net_2931;
wire net_12097;
wire net_6846;
wire net_18250;
wire net_17965;
wire net_598;
wire net_4967;
wire net_18709;
wire net_3455;
wire net_6317;
wire net_12011;
wire net_10068;
wire net_16421;
wire net_18438;
wire net_4818;
wire net_2820;
wire net_8690;
wire net_6091;
wire net_8348;
wire net_18914;
wire net_18689;
wire net_4404;
wire net_3068;
wire net_5973;
wire net_8585;
wire net_3892;
wire net_7921;
wire net_18183;
wire net_7080;
wire net_17911;
wire net_5978;
wire net_6739;
wire net_632;
wire net_843;
wire net_3860;
wire net_15652;
wire net_15603;
wire net_12720;
wire net_16759;
wire net_10063;
wire x661;
wire net_5484;
wire net_2100;
wire net_11959;
wire net_2122;
wire net_6617;
wire net_12572;
wire net_18396;
wire net_1540;
wire net_9734;
wire net_11835;
wire net_18655;
wire net_1725;
wire net_10393;
wire net_3541;
wire net_16532;
wire net_18789;
wire net_5649;
wire net_3532;
wire net_13718;
wire net_12725;
wire net_17307;
wire net_5112;
wire net_18149;
wire net_17700;
wire net_5190;
wire net_9750;
wire net_10303;
wire net_6554;
wire net_14712;
wire net_503;
wire net_7504;
wire net_16676;
wire net_13510;
wire net_18798;
wire net_5695;
wire net_2103;
wire net_1672;
wire net_11818;
wire net_996;
wire net_3091;
wire net_14165;
wire net_2994;
wire net_16510;
wire net_11617;
wire net_10838;
wire net_8327;
wire net_17504;
wire net_4004;
wire net_8767;
wire net_7706;
wire net_18705;
wire net_18605;
wire net_2973;
wire net_9304;
wire net_12342;
wire net_3106;
wire net_13792;
wire net_2503;
wire net_16683;
wire net_9705;
wire net_15170;
wire net_6646;
wire net_17834;
wire net_6469;
wire net_13578;
wire net_18565;
wire net_8330;
wire net_9821;
wire net_18889;
wire net_6211;
wire net_13670;
wire net_3721;
wire net_4606;
wire net_10556;
wire net_10982;
wire net_8894;
wire net_6572;
wire net_12397;
wire net_7416;
wire net_11677;
wire net_15064;
wire net_6901;
wire net_14726;
wire net_5051;
wire net_10688;
wire net_2469;
wire net_11214;
wire net_17229;
wire net_14819;
wire net_15938;
wire net_18545;
wire net_17421;
wire net_1404;
wire net_1012;
wire net_10458;
wire net_14824;
wire x4049;
wire net_5807;
wire net_8809;
wire net_4694;
wire net_2036;
wire net_395;
wire net_15124;
wire net_12988;
wire net_15448;
wire net_8070;
wire net_9182;
wire net_10219;
wire net_17064;
wire net_8623;
wire net_2323;
wire net_3867;
wire net_16223;
wire net_3677;
wire net_4811;
wire net_15088;
wire net_16864;
wire net_5451;
wire net_15336;
wire net_4972;
wire net_10599;
wire net_10459;
wire x890;
wire net_17032;
wire net_1901;
wire net_4890;
wire net_8429;
wire net_3021;
wire net_3711;
wire net_7580;
wire net_602;
wire net_4580;
wire net_12605;
wire net_2379;
wire net_8273;
wire net_2918;
wire net_10932;
wire net_12288;
wire net_16084;
wire net_1497;
wire net_11658;
wire net_1800;
wire net_18590;
wire net_4634;
wire net_14480;
wire net_279;
wire net_3347;
wire net_12281;
wire net_18440;
wire net_4039;
wire net_4030;
wire net_11326;
wire net_10212;
wire net_6337;
wire net_10713;
wire net_15506;
wire net_14119;
wire net_4078;
wire net_14289;
wire net_2833;
wire net_2561;
wire net_12170;
wire net_15224;
wire net_17801;
wire net_18326;
wire x13761;
wire net_18007;
wire net_13775;
wire net_17183;
wire net_3813;
wire net_16599;
wire net_18587;
wire net_1531;
wire net_1159;
wire net_10666;
wire net_861;
wire net_10334;
wire net_6755;
wire net_7217;
wire net_12645;
wire net_6696;
wire net_12400;
wire net_11102;
wire net_4914;
wire net_17658;
wire net_8544;
wire net_10882;
wire net_15814;
wire net_5213;
wire net_12951;
wire net_7696;
wire net_8567;
wire net_4552;
wire net_16946;
wire net_1527;
wire net_18963;
wire net_13270;
wire net_268;
wire net_11849;
wire net_3386;
wire net_4134;
wire net_6631;
wire net_13324;
wire net_15627;
wire net_9406;
wire net_17135;
wire net_17117;
wire net_14536;
wire net_3638;
wire net_2570;
wire net_19040;
wire net_5793;
wire net_3354;
wire net_13195;
wire net_16558;
wire net_9468;
wire net_2712;
wire net_2005;
wire net_13976;
wire net_14827;
wire net_2771;
wire net_1123;
wire net_4897;
wire net_6040;
wire net_18947;
wire net_9343;
wire net_13911;
wire net_9980;
wire net_11241;
wire net_4838;
wire net_5958;
wire net_3363;
wire net_984;
wire net_11894;
wire net_5467;
wire net_6407;
wire net_7263;
wire net_10915;
wire net_13652;
wire net_1105;
wire net_12370;
wire net_2172;
wire net_11448;
wire net_14023;
wire net_15904;
wire net_16718;
wire net_7491;
wire net_18407;
wire net_4457;
wire net_9519;
wire net_1856;
wire net_830;
wire net_16205;
wire net_1279;
wire net_14642;
wire net_1047;
wire net_18019;
wire net_13003;
wire net_9475;
wire net_18523;
wire net_18080;
wire net_12642;
wire net_6394;
wire net_8439;
wire net_18698;
wire net_14553;
wire net_4688;
wire net_11425;
wire net_17339;
wire net_2631;
wire net_8101;
wire net_16129;
wire net_16906;
wire net_12386;
wire net_12926;
wire net_1467;
wire net_3181;
wire net_1061;
wire net_5623;
wire net_5951;
wire net_18121;
wire net_3837;
wire net_9096;
wire net_2288;
wire net_4839;
wire net_14843;
wire net_8718;
wire net_13752;
wire net_11189;
wire net_15213;
wire net_18763;
wire net_17414;
wire net_16320;
wire net_17681;
wire net_15200;
wire net_3983;
wire net_14378;
wire net_8121;
wire net_3814;
wire net_15730;
wire net_10534;
wire net_6266;
wire net_2072;
wire net_18691;
wire net_1872;
wire net_16233;
wire net_1716;
wire net_13926;
wire net_5003;
wire net_1607;
wire net_5247;
wire net_11768;
wire net_13472;
wire net_17222;
wire net_1263;
wire net_16377;
wire net_12331;
wire net_17924;
wire net_3452;
wire net_196;
wire net_4591;
wire net_8766;
wire net_11969;
wire net_14356;
wire net_2067;
wire net_8120;
wire net_14243;
wire net_8881;
wire net_5183;
wire net_7200;
wire net_18098;
wire net_1639;
wire net_16193;
wire net_5267;
wire net_4126;
wire net_4549;
wire net_7284;
wire net_3625;
wire net_11431;
wire net_14435;
wire net_4145;
wire net_7604;
wire x13115;
wire net_15145;
wire net_2152;
wire net_732;
wire net_11981;
wire net_12880;
wire net_5286;
wire net_6105;
wire net_8285;
wire net_2088;
wire net_13083;
wire net_6423;
wire net_7572;
wire net_13963;
wire net_2689;
wire net_4217;
wire net_10655;
wire net_17646;
wire net_17121;
wire net_8422;
wire net_11678;
wire net_15399;
wire net_11092;
wire x12891;
wire net_15935;
wire net_13970;
wire net_449;
wire net_5234;
wire net_8225;
wire net_11523;
wire net_1087;
wire net_15697;
wire net_18806;
wire net_4234;
wire net_11064;
wire net_3995;
wire net_733;
wire net_887;
wire net_8245;
wire net_5856;
wire net_18011;
wire net_18865;
wire x3524;
wire net_6098;
wire net_7537;
wire net_11975;
wire net_6151;
wire net_10491;
wire net_2308;
wire net_6301;
wire net_9105;
wire net_4628;
wire net_2770;
wire net_2636;
wire net_1424;
wire net_4375;
wire net_19043;
wire net_4412;
wire net_16840;
wire net_9287;
wire net_17391;
wire net_18834;
wire net_8167;
wire net_4280;
wire net_10347;
wire net_9563;
wire net_950;
wire x240;
wire net_11441;
wire x338;
wire net_9839;
wire net_2816;
wire net_17435;
wire net_6610;
wire net_7651;
wire net_14507;
wire net_18959;
wire net_14344;
wire net_1214;
wire net_3641;
wire net_9529;
wire net_866;
wire net_12895;
wire net_4220;
wire net_12700;
wire net_15705;
wire net_10681;
wire net_18704;
wire net_18047;
wire net_1032;
wire net_567;
wire net_15563;
wire net_13985;
wire net_3726;
wire net_5255;
wire net_18506;
wire net_272;
wire net_5787;
wire net_13345;
wire net_8458;
wire net_13384;
wire net_3939;
wire net_14625;
wire net_1024;
wire net_12480;
wire net_1590;
wire x13093;
wire net_14097;
wire net_18495;
wire net_1612;
wire net_17268;
wire net_814;
wire net_11121;
wire net_13685;
wire net_17320;
wire x13733;
wire net_5840;
wire net_8128;
wire net_6184;
wire net_12705;
wire net_12525;
wire net_17641;
wire net_14003;
wire net_3930;
wire net_4785;
wire net_10639;
wire net_9815;
wire net_3299;
wire net_2586;
wire net_15795;
wire net_1655;
wire net_10290;
wire net_6963;
wire net_2365;
wire net_15951;
wire net_17803;
wire net_18306;
wire net_17179;
wire net_4797;
wire net_9240;
wire net_10810;
wire net_2598;
wire net_2361;
wire net_18031;
wire net_11194;
wire net_14767;
wire net_17717;
wire net_2879;
wire net_1680;
wire net_14219;
wire net_16172;
wire net_16258;
wire net_3302;
wire net_17481;
wire net_7540;
wire net_15276;
wire net_15925;
wire net_11337;
wire net_3187;
wire net_15250;
wire net_2622;
wire net_5966;
wire net_10514;
wire net_8294;
wire net_17690;
wire net_10997;
wire net_14500;
wire net_2262;
wire net_7505;
wire net_2087;
wire net_1002;
wire net_7620;
wire net_7224;
wire net_6118;
wire net_3188;
wire net_13308;
wire net_17259;
wire net_1993;
wire net_8198;
wire x2195;
wire net_11128;
wire net_8724;
wire net_2903;
wire net_8683;
wire net_11623;
wire net_8392;
wire net_9556;
wire net_4128;
wire net_16262;
wire net_4923;
wire net_3873;
wire net_11866;
wire net_6015;
wire net_2155;
wire net_6741;
wire net_168;
wire net_15056;
wire net_17194;
wire net_385;
wire net_2609;
wire net_13253;
wire net_14179;
wire net_5365;
wire net_5736;
wire net_5404;
wire net_5044;
wire net_14890;
wire net_8657;
wire net_10260;
wire net_8139;
wire x4821;
wire net_10468;
wire net_6236;
wire net_11220;
wire net_7660;
wire net_13675;
wire net_2380;
wire net_3393;
wire net_4548;
wire net_8231;
wire net_16031;
wire net_9323;
wire net_16135;
wire net_14797;
wire net_1412;
wire net_16524;
wire net_17816;
wire net_15402;
wire net_12327;
wire net_12965;
wire net_13357;
wire net_7358;
wire net_7211;
wire net_16666;
wire net_3040;
wire net_3557;
wire net_10825;
wire net_13762;
wire net_10609;
wire net_15975;
wire net_8801;
wire net_3004;
wire net_18453;
wire net_8014;
wire net_12624;
wire net_7244;
wire net_17631;
wire net_7981;
wire net_10315;
wire net_16500;
wire net_3830;
wire net_9757;
wire net_8464;
wire net_17756;
wire net_12561;
wire net_12806;
wire net_10282;
wire net_18177;
wire net_833;
wire net_14044;
wire net_12744;
wire net_6656;
wire net_17914;
wire net_4758;
wire net_4249;
wire net_14512;
wire net_14757;
wire net_12931;
wire net_1399;
wire net_11349;
wire net_13681;
wire net_16270;
wire net_8529;
wire net_8667;
wire net_3350;
wire net_15877;
wire net_3553;
wire net_5161;
wire net_14489;
wire net_16578;
wire net_7623;
wire net_15416;
wire net_16277;
wire net_12751;
wire net_1781;
wire net_16067;
wire x13950;
wire net_18998;
wire net_3049;
wire net_7457;
wire net_10299;
wire net_6918;
wire net_17572;
wire net_2514;
wire net_9250;
wire net_12183;
wire net_3474;
wire net_4775;
wire net_16754;
wire net_2013;
wire net_5472;
wire net_15990;
wire net_7477;
wire net_13503;
wire net_11262;
wire net_18556;
wire net_17869;
wire net_2028;
wire net_9758;
wire net_1889;
wire net_3766;
wire net_7361;
wire net_12065;
wire net_8717;
wire net_2981;
wire net_17895;
wire net_1164;
wire net_6810;
wire net_8912;
wire net_10817;
wire net_15528;
wire x4757;
wire net_14449;
wire net_6923;
wire net_11148;
wire net_12500;
wire net_2583;
wire x4667;
wire net_5708;
wire net_8854;
wire net_4665;
wire net_5824;
wire net_9366;
wire net_16525;
wire net_2706;
wire net_5163;
wire net_5580;
wire net_11842;
wire net_8304;
wire net_2602;
wire net_6366;
wire net_8449;
wire net_17970;
wire net_4484;
wire net_440;
wire net_8069;
wire net_8048;
wire net_10866;
wire net_17021;
wire net_5664;
wire net_14747;
wire net_16799;
wire net_4652;
wire net_14558;
wire net_718;
wire net_6178;
wire net_7773;
wire net_18023;
wire net_18243;
wire net_14193;
wire net_8707;
wire net_5714;
wire net_12995;
wire net_13367;
wire net_5838;
wire net_12215;
wire net_13946;
wire net_17579;
wire x132;
wire net_13545;
wire net_14078;
wire net_4448;
wire net_16985;
wire net_336;
wire net_9419;
wire net_15598;
wire net_10404;
wire net_14033;
wire net_1578;
wire net_14584;
wire net_18464;
wire x13843;
wire net_8417;
wire net_18206;
wire net_17097;
wire net_697;
wire net_2003;
wire net_5053;
wire net_18288;
wire net_17410;
wire net_3426;
wire net_13008;
wire net_15632;
wire net_5095;
wire net_1333;
wire net_5325;
wire net_5924;
wire net_18483;
wire net_5107;
wire net_5593;
wire net_17662;
wire net_3082;
wire net_14422;
wire net_5859;
wire net_10802;
wire net_11503;
wire net_3676;
wire net_13521;
wire net_4185;
wire net_4204;
wire net_5630;
wire net_6072;
wire net_7591;
wire net_2054;
wire net_6682;
wire net_9880;
wire net_17665;
wire net_6295;
wire net_9133;
wire net_14057;
wire net_10901;
wire net_14133;
wire net_15160;
wire net_2793;
wire net_18459;
wire net_1836;
wire net_14971;
wire net_4310;
wire net_8783;
wire net_10570;
wire net_5922;
wire net_13158;
wire net_14571;
wire net_3430;
wire net_11557;
wire net_8266;
wire net_6795;
wire net_15016;
wire net_4244;
wire net_14882;
wire net_18220;
wire net_7887;
wire net_15779;
wire net_6930;
wire net_4396;
wire net_6158;
wire net_9273;
wire net_16361;
wire net_2398;
wire net_4581;
wire net_7811;
wire net_12140;
wire x13374;
wire net_4431;
wire net_7821;
wire net_15374;
wire net_3315;
wire net_16580;
wire net_2455;
wire net_17624;
wire net_12732;
wire net_17400;
wire net_10753;
wire net_8493;
wire net_8744;
wire net_18124;
wire net_1386;
wire net_7841;
wire net_9431;
wire net_6546;
wire net_8949;
wire net_6115;
wire net_16150;
wire net_10550;
wire net_12805;
wire net_5991;
wire net_5101;
wire net_10252;
wire net_14968;
wire net_14989;
wire net_2186;
wire net_3696;
wire net_3473;
wire net_13551;
wire net_17231;
wire net_569;
wire net_12062;
wire net_13877;
wire net_16781;
wire net_12767;
wire net_8857;
wire x4496;
wire net_4018;
wire net_17439;
wire net_17281;
wire net_6826;
wire net_15249;
wire net_13696;
wire net_18710;
wire net_3124;
wire net_1903;
wire net_2407;
wire net_13467;
wire net_10600;
wire net_13162;
wire net_7412;
wire net_13414;
wire net_17907;
wire net_2078;
wire net_779;
wire net_16511;
wire net_12473;
wire net_14438;
wire net_234;
wire net_4151;
wire net_12634;
wire net_5142;
wire net_13258;
wire net_17126;
wire net_16632;
wire net_15309;
wire net_5764;
wire net_7390;
wire net_11469;
wire net_17653;
wire net_7732;
wire net_6583;
wire net_9128;
wire net_491;
wire net_11460;
wire net_1299;
wire net_948;
wire net_6679;
wire net_18599;
wire net_11573;
wire net_17462;
wire net_17109;
wire net_2593;
wire net_876;
wire net_6479;
wire net_15841;
wire net_2162;
wire net_18820;
wire net_10833;
wire net_15424;
wire net_7154;
wire net_9646;
wire net_16041;
wire net_8601;
wire net_11960;
wire net_1458;
wire net_18160;
wire net_5587;
wire net_17160;
wire net_10184;
wire net_5933;
wire net_16977;
wire net_905;
wire net_10591;
wire net_14122;
wire net_2229;
wire net_158;
wire net_5774;
wire net_10613;
wire net_13842;
wire net_7370;
wire net_3200;
wire net_14848;
wire net_19039;
wire net_16181;
wire net_15457;
wire net_5624;
wire net_16011;
wire net_2504;
wire net_11571;
wire net_2175;
wire net_3784;
wire net_5650;
wire net_18882;
wire net_10214;
wire net_15637;
wire net_2116;
wire net_4327;
wire net_14701;
wire net_11334;
wire net_8035;
wire net_16973;
wire net_8090;
wire net_9572;
wire net_1967;
wire net_11565;
wire net_5171;
wire net_9333;
wire net_6860;
wire net_8754;
wire net_16481;
wire net_465;
wire net_14676;
wire net_1883;
wire net_17948;
wire net_11233;
wire net_17381;
wire net_3058;
wire net_8484;
wire net_1315;
wire net_6994;
wire net_5904;
wire net_5358;
wire net_10073;
wire net_15790;
wire net_5208;
wire net_9767;
wire net_5019;
wire net_13144;
wire net_6956;
wire net_9376;
wire net_9903;
wire x13156;
wire net_4977;
wire net_10138;
wire net_5075;
wire net_11646;
wire net_7327;
wire net_293;
wire net_15117;
wire net_3666;
wire net_11890;
wire net_1938;
wire net_13303;
wire net_15677;
wire net_1823;
wire net_14660;
wire net_5081;
wire net_15516;
wire net_3576;
wire net_191;
wire net_558;
wire net_2069;
wire net_15021;
wire net_1618;
wire net_10910;
wire net_14399;
wire net_2497;
wire net_11594;
wire net_3562;
wire net_7006;
wire net_15319;
wire net_15110;
wire net_5885;
wire net_7112;
wire net_11905;
wire net_18893;
wire net_4023;
wire net_14720;
wire net_15853;
wire net_7755;
wire net_4450;
wire net_6881;
wire net_15610;
wire net_6942;
wire net_1984;
wire net_13959;
wire net_4670;
wire net_10734;
wire net_16436;
wire net_1944;
wire net_11545;
wire net_1775;
wire net_10112;
wire net_16993;
wire net_297;
wire net_346;
wire net_10158;
wire net_17956;
wire net_10693;
wire net_13725;
wire net_15982;
wire net_15870;
wire net_229;
wire net_14835;
wire net_4360;
wire net_4962;
wire net_687;
wire x4347;
wire net_17334;
wire net_15073;
wire net_3266;
wire net_4160;
wire net_13339;
wire net_14702;
wire net_17265;
wire net_3888;
wire net_7072;
wire net_13949;
wire net_14303;
wire net_3566;
wire net_15263;
wire net_14945;
wire net_3596;
wire net_10143;
wire net_5021;
wire net_13741;
wire net_9296;
wire net_9345;
wire net_5415;
wire net_1184;
wire net_13492;
wire net_4055;
wire net_5339;
wire net_18268;
wire net_6482;
wire net_18924;
wire net_6961;
wire net_14444;
wire net_7383;
wire net_15363;
wire net_10722;
wire net_5425;
wire net_1960;
wire net_9660;
wire net_15622;
wire net_7435;
wire net_12548;
wire x12955;
wire net_15194;
wire net_828;
wire net_4256;
wire net_9145;
wire net_6222;
wire net_1603;
wire net_4490;
wire net_12222;
wire net_14349;
wire x275;
wire net_13031;
wire net_18728;
wire net_7446;
wire net_10009;
wire net_10108;
wire x577;
wire net_11017;
wire net_18981;
wire net_18321;
wire net_8385;
wire net_3521;
wire net_14877;
wire net_982;
wire net_14874;
wire net_9610;
wire net_1580;
wire net_3896;
wire net_5287;
wire net_4384;
wire net_6462;
wire net_9189;
wire net_17189;
wire net_9314;
wire net_9576;
wire net_4912;
wire net_6002;
wire net_14501;
wire net_15863;
wire net_5748;
wire net_12076;
wire net_15531;
wire net_8180;
wire net_5049;
wire net_10869;
wire net_11393;
wire net_17537;
wire net_11058;
wire net_8899;
wire net_225;
wire net_14927;
wire net_3128;
wire net_4733;
wire net_12937;
wire net_6524;
wire net_5313;
wire net_15334;
wire net_2611;
wire net_871;
wire net_11804;
wire net_14974;
wire net_390;
wire net_1154;
wire net_11789;
wire net_6983;
wire net_6593;
wire net_11782;
wire net_16249;
wire net_4294;
wire net_5128;
wire net_6062;
wire net_15723;
wire net_12735;
wire net_7494;
wire net_12798;
wire net_280;
wire net_12132;
wire net_12027;
wire net_12715;
wire x2100;
wire net_495;
wire net_13022;
wire net_16317;
wire net_10569;
wire net_2140;
wire net_13180;
wire net_6345;
wire net_13975;
wire net_15965;
wire net_16124;
wire net_13211;
wire net_2517;
wire net_8798;
wire net_2316;
wire net_12105;
wire net_8644;
wire net_6457;
wire net_14525;
wire net_6100;
wire net_6356;
wire net_2703;
wire net_11273;
wire net_13524;
wire net_14214;
wire net_1441;
wire net_18814;
wire net_969;
wire net_9154;
wire net_1525;
wire net_7097;
wire net_12710;
wire net_17443;
wire net_11458;
wire net_821;
wire net_4003;
wire net_13444;
wire net_4177;
wire net_9350;
wire net_18302;
wire net_8936;
wire net_8345;
wire net_2335;
wire net_11210;
wire net_3940;
wire net_14603;
wire net_18352;
wire net_11533;
wire net_11161;
wire net_14153;
wire net_2618;
wire net_4316;
wire net_6045;
wire net_6540;
wire net_14688;
wire net_16571;
wire net_7952;
wire net_16497;
wire net_12786;
wire net_8670;
wire net_5411;
wire net_12691;
wire net_1748;
wire net_3078;
wire net_2964;
wire net_11882;
wire net_9946;
wire net_16589;
wire net_2343;
wire net_2232;
wire net_726;
wire net_13241;
wire net_15349;
wire net_3237;
wire net_701;
wire net_808;
wire net_5553;
wire net_9121;
wire net_1704;
wire net_4821;
wire net_5026;
wire net_2738;
wire net_16432;
wire net_2944;
wire net_18624;
wire net_18259;
wire net_12079;
wire net_14384;
wire net_17709;
wire net_6662;
wire net_11176;
wire net_18417;
wire net_9451;
wire net_13058;
wire net_7927;
wire net_17247;
wire net_5654;
wire net_16845;
wire net_13034;
wire net_935;
wire net_8827;
wire net_3116;
wire net_1511;
wire net_645;
wire net_11436;
wire net_14649;
wire net_4071;
wire net_17005;
wire net_14242;
wire net_8825;
wire net_10862;
wire net_17428;
wire net_4533;
wire net_17963;
wire net_17145;
wire net_1816;
wire net_8076;
wire net_4195;
wire net_7909;
wire net_16149;
wire net_14085;
wire net_331;
wire net_12597;
wire net_17853;
wire net_4644;
wire net_8633;
wire net_2220;
wire net_4762;
wire net_2823;
wire net_3728;
wire net_5724;
wire net_7138;
wire net_4884;
wire net_12981;
wire net_8000;
wire net_15537;
wire net_12541;
wire net_15764;
wire net_13808;
wire net_16399;
wire net_12841;
wire net_14333;
wire net_16615;
wire net_12199;
wire net_16928;
wire net_1259;
wire net_4753;
wire net_11207;
wire net_2839;
wire net_2143;
wire net_4225;
wire net_2196;
wire net_3791;
wire net_7676;
wire net_8059;
wire net_10478;
wire net_5275;
wire net_11611;
wire net_478;
wire net_16672;
wire net_6608;
wire net_11429;
wire net_4959;
wire net_5781;
wire net_8733;
wire net_1975;
wire net_8958;
wire net_8375;
wire net_13067;
wire net_11948;
wire net_13991;
wire net_5600;
wire net_17986;
wire net_7406;
wire net_17369;
wire net_7530;
wire net_7253;
wire net_3028;
wire net_18432;
wire net_17073;
wire net_11281;
wire net_1692;
wire net_7087;
wire net_5079;
wire net_12675;
wire net_2655;
wire net_2528;
wire net_16588;
wire net_18100;
wire net_10854;
wire net_9682;
wire net_1361;
wire net_16744;
wire net_2450;
wire net_9260;
wire net_14118;
wire net_1208;
wire net_7948;
wire net_16161;
wire net_8920;
wire net_13201;
wire net_12162;
wire net_18600;
wire x13077;
wire net_8560;
wire net_13769;
wire net_9279;
wire net_12954;
wire net_4710;
wire net_13378;
wire net_18780;
wire net_4808;
wire net_13810;
wire net_2889;
wire net_5506;
wire net_9537;
wire net_16731;
wire net_4544;
wire net_17887;
wire net_16504;
wire net_7340;
wire net_13901;
wire net_12187;
wire net_6398;
wire net_3154;
wire net_4828;
wire net_15568;
wire net_15929;
wire net_16088;
wire net_9862;
wire net_3622;
wire net_13190;
wire net_9800;
wire net_10398;
wire net_2729;
wire net_10389;
wire net_4422;
wire net_16251;
wire net_10116;
wire net_302;
wire net_18954;
wire net_1131;
wire net_753;
wire net_17283;
wire net_15668;
wire net_9034;
wire net_5575;
wire net_18330;
wire net_9710;
wire x4778;
wire net_12464;
wire net_13609;
wire net_8084;
wire net_4155;
wire net_13864;
wire net_6353;
wire net_11297;
wire x4576;
wire net_6722;
wire net_8288;
wire net_6283;
wire net_12861;
wire net_5192;
wire net_12301;
wire net_13268;
wire net_1228;
wire net_10146;
wire net_7148;
wire net_17386;
wire net_7807;
wire net_2722;
wire net_13092;
wire net_16455;
wire net_9891;
wire net_12139;
wire net_6504;
wire net_9399;
wire net_8531;
wire net_12013;
wire net_13113;
wire net_16419;
wire net_15190;
wire net_8536;
wire net_11548;
wire net_11380;
wire net_17858;
wire net_13602;
wire net_11795;
wire net_1057;
wire net_2915;
wire net_17808;
wire net_7235;
wire net_15673;
wire net_5225;
wire net_10895;
wire net_6161;
wire net_6953;
wire net_2987;
wire net_10647;
wire net_15199;
wire net_18759;
wire net_2253;
wire net_1699;
wire net_9534;
wire net_4792;
wire net_12944;
wire net_13267;
wire net_15589;
wire net_11133;
wire net_11309;
wire net_16959;
wire net_18649;
wire net_2521;
wire net_6246;
wire net_12915;
wire net_11296;
wire net_1016;
wire net_16410;
wire net_6437;
wire net_9035;
wire net_15256;
wire net_10017;
wire net_11315;
wire net_16970;
wire net_18248;
wire net_3977;
wire net_10323;
wire net_4567;
wire x1070;
wire net_1744;
wire net_10201;
wire net_10417;
wire net_18664;
wire net_516;
wire net_17532;
wire net_3176;
wire net_3585;
wire net_11776;
wire net_12655;
wire net_12614;
wire net_956;
wire net_3963;
wire net_5799;
wire net_14383;
wire net_5496;
wire net_438;
wire net_15770;
wire net_8181;
wire net_18062;
wire net_8178;
wire net_18668;
wire net_2250;
wire net_12334;
wire net_3013;
wire net_5278;
wire net_5438;
wire net_13826;
wire net_3110;
wire net_2967;
wire net_10916;
wire net_8214;
wire net_13337;
wire net_17020;
wire net_7598;
wire net_6808;
wire net_18227;
wire net_10645;
wire net_13185;
wire net_17360;
wire net_15471;
wire net_3570;
wire net_15283;
wire net_17081;
wire x815;
wire net_15663;
wire net_15678;
wire net_5916;
wire net_9773;
wire net_18991;
wire net_2785;
wire net_9693;
wire net_10840;
wire net_8575;
wire net_473;
wire net_8274;
wire net_13169;
wire net_18467;
wire net_18745;
wire net_3599;
wire net_14426;
wire net_16012;
wire net_5099;
wire net_8350;
wire net_9512;
wire x352;
wire net_454;
wire net_5349;
wire net_6251;
wire net_15518;
wire net_16384;
wire net_18036;
wire net_709;
wire net_2484;
wire net_13535;
wire net_11342;
wire net_10791;
wire net_1066;
wire net_5514;
wire net_9956;
wire net_15095;
wire net_4304;
wire net_5847;
wire net_1344;
wire net_4560;
wire net_1084;
wire net_1500;
wire net_9778;
wire net_1136;
wire net_11376;
wire net_5418;
wire net_14010;
wire net_3008;
wire net_2763;
wire net_11707;
wire net_573;
wire net_18277;
wire net_9065;
wire net_12412;
wire net_6855;
wire net_13314;
wire net_15912;
wire net_17069;
wire net_3616;
wire net_11606;
wire net_9494;
wire net_17677;
wire net_5521;
wire net_8570;
wire net_13352;
wire net_5037;
wire net_3672;
wire net_6089;
wire net_11101;
wire net_9249;
wire net_14371;
wire net_11879;
wire net_5811;
wire net_941;
wire net_7560;
wire net_6038;
wire net_13292;
wire net_14351;
wire net_14582;
wire net_8129;
wire net_2311;
wire net_17054;
wire net_9444;
wire net_4611;
wire net_7500;
wire net_17214;
wire net_1599;
wire net_6587;
wire net_10575;
wire net_15151;
wire net_11087;
wire net_17242;
wire net_3828;
wire net_3132;
wire net_11504;
wire net_9973;
wire net_12240;
wire net_3053;
wire net_9802;
wire net_15209;
wire net_9579;
wire net_7187;
wire net_7460;
wire net_6601;
wire net_2023;
wire net_8518;
wire net_4523;
wire net_13923;
wire net_15041;
wire net_262;
wire net_527;
wire net_1668;
wire net_12151;
wire net_7552;
wire net_3139;
wire net_4063;
wire net_5388;
wire net_6399;
wire net_16362;
wire net_1793;
wire net_11714;
wire net_18092;
wire net_3786;
wire net_7161;
wire net_8261;
wire net_6215;
wire net_5706;
wire net_1859;
wire net_145;
wire net_12550;
wire net_15299;
wire net_8193;
wire net_10699;
wire net_10431;
wire net_2804;
wire net_4637;
wire net_11134;
wire net_188;
wire net_5535;
wire net_3753;
wire net_17699;
wire net_3319;
wire net_4353;
wire net_18855;
wire net_16425;
wire net_10160;
wire net_7141;
wire net_1077;
wire net_2924;
wire net_6520;
wire net_14163;
wire net_8969;
wire net_10050;
wire net_15700;
wire net_17638;
wire net_12318;
wire net_8022;
wire net_11825;
wire net_2410;
wire net_8281;
wire net_16913;
wire net_9208;
wire net_3108;
wire net_18423;
wire net_16895;
wire net_10975;
wire net_2185;
wire net_10445;
wire net_13103;
wire net_1321;
wire net_15780;
wire net_14263;
wire net_4441;
wire x378;
wire net_5392;
wire net_8741;
wire net_4949;
wire net_14484;
wire net_1099;
wire net_18384;
wire net_7106;
wire net_14901;
wire net_17378;
wire net_7103;
wire net_14543;
wire net_9227;
wire net_9885;
wire net_18586;
wire net_404;
wire net_15185;
wire net_11683;
wire net_6033;
wire net_14941;
wire net_5455;
wire net_11624;
wire net_2666;
wire net_9276;
wire net_10929;
wire net_8402;
wire net_18715;
wire net_1239;
wire net_8663;
wire net_10246;
wire net_1463;
wire net_9743;
wire net_8793;
wire net_12257;
wire net_17825;
wire net_15833;
wire net_10081;
wire net_9266;
wire net_17325;
wire net_3822;
wire net_15139;
wire x4115;
wire net_17015;
wire net_6872;
wire net_16054;
wire net_484;
wire net_896;
wire net_18156;
wire net_7655;
wire net_3223;
wire net_5894;
wire net_11363;
wire net_11599;
wire net_16960;
wire net_15135;
wire net_10088;
wire net_9795;
wire net_18547;
wire net_12971;
wire net_13106;
wire net_11563;
wire net_11794;
wire net_13939;
wire net_15031;
wire net_7917;
wire net_11550;
wire net_13614;
wire net_1896;
wire net_1982;
wire net_14577;
wire net_13283;
wire net_12687;
wire net_16604;
wire net_16330;
wire net_8089;
wire net_12084;
wire net_10014;
wire net_15960;
wire net_11719;
wire net_6509;
wire net_12507;
wire net_3253;
wire net_10630;
wire net_6935;
wire net_5498;
wire net_13176;
wire net_1882;
wire net_12347;
wire net_12229;
wire net_12755;
wire net_7744;
wire net_16967;
wire net_413;
wire net_11072;
wire net_9613;
wire net_18540;
wire net_6141;
wire net_14982;
wire net_12666;
wire x1130;
wire net_2419;
wire net_7876;
wire net_10154;
wire net_5753;
wire net_14898;
wire net_7608;
wire net_12203;
wire net_14315;
wire net_18334;
wire net_253;
wire net_276;
wire net_11696;
wire net_9728;
wire net_14229;
wire net_17453;
wire net_8470;
wire net_12112;
wire net_13899;
wire net_15800;
wire net_6490;
wire net_10586;
wire net_16347;
wire net_9799;
wire net_13395;
wire net_616;
wire net_17977;
wire net_18086;
wire net_1847;
wire net_18772;
wire net_17474;
wire net_17270;
wire net_15899;
wire net_2717;
wire net_793;
wire x324;
wire net_9137;
wire net_2353;
wire net_2272;
wire net_11919;
wire net_9231;
wire net_16934;
wire net_9708;
wire net_4104;
wire net_3287;
wire net_8133;
wire net_14922;
wire net_11305;
wire net_16465;
wire net_2866;
wire net_5866;
wire net_17787;
wire net_18651;
wire net_3025;
wire net_5407;
wire net_17568;
wire net_7673;
wire net_7309;
wire net_6071;
wire net_10342;
wire net_17131;
wire net_6894;
wire net_205;
wire net_1286;
wire net_11702;
wire net_6427;
wire net_15204;
wire net_9764;
wire net_11872;
wire net_15290;
wire net_17780;
wire net_7617;
wire net_18955;
wire net_7533;
wire net_1952;
wire net_18497;
wire net_9214;
wire net_9846;
wire net_11495;
wire net_12512;
wire net_4620;
wire net_380;
wire net_5696;
wire net_14141;
wire net_2847;
wire net_6515;
wire net_7932;
wire net_1556;
wire net_12885;
wire net_5911;
wire net_6803;
wire net_4337;
wire net_13548;
wire net_7976;
wire net_16292;
wire net_4745;
wire net_1270;
wire net_17610;
wire net_16657;
wire net_4905;
wire net_15345;
wire net_18613;
wire net_9717;
wire net_14178;
wire net_6094;
wire net_14454;
wire net_18375;
wire net_7712;
wire net_17043;
wire net_3878;
wire net_4940;
wire net_8132;
wire net_5585;
wire net_3241;
wire net_7273;
wire net_17748;
wire net_2555;
wire net_4864;
wire net_3504;
wire net_18490;
wire net_1687;
wire net_16857;
wire net_1762;
wire net_5243;
wire net_7407;
wire net_18910;
wire net_1181;
wire net_10685;
wire net_12299;
wire net_313;
wire net_932;
wire net_7472;
wire net_15577;
wire net_6082;
wire net_16446;
wire net_10783;
wire net_13403;
wire net_12488;
wire net_4767;
wire net_5271;
wire net_14257;
wire net_6771;
wire net_12814;
wire net_972;
wire net_7769;
wire net_17526;
wire net_9650;
wire net_15043;
wire net_4725;
wire net_15942;
wire net_6201;
wire net_11669;
wire net_14292;
wire net_7047;
wire net_1489;
wire net_13665;
wire net_15789;
wire net_4343;
wire net_10276;
wire net_16282;
wire net_7794;
wire net_2392;
wire net_7194;
wire net_17515;
wire net_10278;
wire net_8441;
wire net_13064;
wire net_10266;
wire net_1040;
wire net_5947;
wire net_8978;
wire net_6781;
wire net_3089;
wire net_3037;
wire net_4472;
wire net_4463;
wire net_7331;
wire net_18115;
wire net_3686;
wire net_2907;
wire net_15607;
wire net_2243;
wire net_379;
wire net_1569;
wire net_16951;
wire net_3133;
wire net_7795;
wire net_2559;
wire net_18614;
wire net_14451;
wire net_14475;
wire net_1358;
wire net_8477;
wire net_6815;
wire net_14708;
wire net_11405;
wire net_6888;
wire net_8927;
wire net_8421;
wire net_16409;
wire net_960;
wire net_3704;
wire net_17352;
wire net_8155;
wire net_10706;
wire net_14957;
wire net_11051;
wire net_14062;
wire net_16468;
wire net_12842;
wire net_13365;
wire net_9445;
wire net_13996;
wire net_6441;
wire net_4348;
wire net_4526;
wire net_7832;
wire net_581;
wire net_8991;
wire net_9909;
wire net_10564;
wire net_13967;
wire net_2899;
wire net_8799;
wire net_17881;
wire net_9609;
wire net_12421;
wire net_658;
wire net_18554;
wire net_7978;
wire net_14565;
wire net_13529;
wire net_2090;
wire net_18294;
wire net_16508;
wire x13341;
wire net_7723;
wire net_9540;
wire net_12509;
wire net_18239;
wire x1039;
wire net_12758;
wire net_10259;
wire net_5801;
wire net_7026;
wire net_8999;
wire net_15270;
wire net_5461;
wire net_1176;
wire net_2676;
wire net_14853;
wire net_6372;
wire net_4989;
wire net_7032;
wire net_11609;
wire net_15949;
wire net_1751;
wire net_13593;
wire net_6733;
wire net_16216;
wire net_3508;
wire net_16401;
wire net_2434;
wire net_2032;
wire net_17843;
wire net_2467;
wire net_17741;
wire net_11524;
wire net_14499;
wire net_14415;
wire net_9916;
wire net_12008;
wire net_17496;
wire net_7223;
wire net_8865;
wire net_17871;
wire net_18640;
wire net_246;
wire net_6613;
wire net_11269;
wire net_13041;
wire net_10121;
wire net_13436;
wire net_14914;
wire net_16140;
wire net_17347;
wire net_6725;
wire net_8968;
wire net_1378;
wire net_1600;
wire net_2531;
wire net_16339;
wire net_12440;
wire net_17720;
wire net_11971;
wire net_15743;
wire net_676;
wire net_11254;
wire net_12492;
wire net_6626;
wire net_4263;
wire net_15592;
wire net_2538;
wire net_17710;
wire net_5133;
wire net_5542;
wire net_5370;
wire net_4260;
wire net_3492;
wire net_2462;
wire net_6010;
wire net_12760;
wire net_9018;
wire net_9635;
wire net_8820;
wire net_3324;
wire net_13485;
wire net_18166;
wire net_16773;
wire net_5426;
wire net_6450;
wire net_6138;
wire net_6979;
wire net_8398;
wire net_7893;
wire net_9600;
wire net_14463;
wire net_8112;
wire net_10429;
wire net_7939;
wire net_11274;
wire net_3207;
wire net_7810;
wire net_13920;
wire net_2204;
wire net_9668;
wire net_5088;
wire net_2492;
wire net_15485;
wire net_9088;
wire net_11188;
wire net_16871;
wire net_16727;
wire net_4045;
wire net_3843;
wire net_15228;
wire net_10223;
wire x1032;
wire net_16048;
wire net_6543;
wire net_7635;
wire net_11005;
wire net_3038;
wire net_2690;
wire net_13560;
wire net_3924;
wire net_7016;
wire net_9825;
wire net_5226;
wire net_10230;
wire net_8811;
wire net_1051;
wire net_10546;
wire net_18984;
wire net_10048;
wire net_10386;
wire net_14770;
wire net_7644;
wire net_7858;
wire net_11034;
wire net_1515;
wire net_1573;
wire net_7669;
wire net_10356;
wire net_18844;
wire net_4983;
wire net_6869;
wire net_13932;
wire net_9984;
wire net_305;
wire net_7100;
wire net_4208;
wire net_4515;
wire net_12433;
wire net_12016;
wire net_15434;
wire net_12452;
wire net_9166;
wire net_16833;
wire net_1125;
wire net_14716;
wire net_18872;
wire net_10195;
wire net_15084;
wire net_10667;
wire net_17236;
wire net_17686;
wire net_12405;
wire net_6687;
wire net_8818;
wire net_15555;
wire net_13592;
wire net_17254;
wire net_18356;
wire net_9175;
wire net_3485;
wire x13541;
wire net_17483;
wire net_16168;
wire net_2886;
wire net_14408;
wire net_1921;
wire net_10945;
wire net_3853;
wire net_16472;
wire net_9962;
wire net_14781;
wire net_15462;
wire net_2135;
wire net_9091;
wire net_667;
wire net_18413;
wire net_853;
wire net_212;
wire x3485;
wire net_12265;
wire net_914;
wire net_9508;
wire net_10254;
wire net_9923;
wire net_12835;
wire net_6320;
wire net_15245;
wire net_6448;
wire x2400;
wire net_875;
wire net_17942;
wire net_5619;
wire net_14807;
wire net_1092;
wire net_627;
wire net_18937;
wire net_18570;
wire net_8759;
wire net_16115;
wire net_15313;
wire net_18388;
wire net_17358;
wire net_15989;
wire net_11042;
wire net_15444;
wire x3156;
wire net_5636;
wire net_15469;
wire net_2473;
wire net_12231;
wire net_16034;
wire net_399;
wire net_8107;
wire net_15284;
wire net_5949;
wire net_5069;
wire net_1390;
wire net_10678;
wire net_5565;
wire net_7180;
wire net_16805;
wire net_10517;
wire net_1112;
wire x1016;
wire net_10747;
wire net_15483;
wire net_5449;
wire net_8146;
wire net_11200;
wire net_12085;
wire net_18191;
wire net_3230;
wire net_13295;
wire net_14494;
wire net_10187;
wire net_8316;
wire net_13585;
wire net_14932;
wire net_5677;
wire net_11486;
wire net_17154;
wire net_5296;
wire net_1310;
wire net_14171;
wire net_9634;
wire net_6057;
wire net_15687;
wire net_18674;
wire net_1304;
wire net_7579;
wire net_4381;
wire net_9471;
wire net_6674;
wire net_11378;
wire net_11918;
wire net_7863;
wire net_13427;
wire net_11450;
wire net_11587;
wire net_10370;
wire net_6127;
wire net_6058;
wire x13626;
wire net_13417;
wire net_10919;
wire net_6070;
wire net_2449;
wire net_17105;
wire net_6588;
wire net_416;
wire net_15986;
wire net_5629;
wire net_16326;
wire net_6896;
wire net_15851;
wire net_6642;
wire net_14814;
wire net_10760;
wire net_1786;
wire net_1377;
wire net_5620;
wire net_16239;
wire net_10253;
wire net_12031;
wire net_4513;
wire net_10940;
wire net_14025;
wire net_5965;
wire net_14439;
wire net_5586;
wire net_11118;
wire net_13428;
wire net_5430;
wire net_17903;
wire net_1393;
wire net_13724;
wire net_17994;
wire net_2169;
wire net_1324;
wire net_8758;
wire net_7114;
wire net_12058;
wire net_8017;
wire net_6997;
wire net_4323;
wire net_9336;
wire net_3527;
wire net_1138;
wire net_8805;
wire net_17598;
wire net_10167;
wire net_18621;
wire x3028;
wire net_3292;
wire net_1439;
wire net_8714;
wire net_13489;
wire net_1778;
wire net_508;
wire net_9700;
wire net_15428;
wire net_6907;
wire net_5098;
wire net_7438;
wire net_15617;
wire net_5355;
wire net_8149;
wire net_11453;
wire net_11962;
wire net_5413;
wire net_4434;
wire net_18128;
wire net_12068;
wire net_16197;
wire net_4744;
wire net_18178;
wire net_6636;
wire net_2896;
wire net_14707;
wire net_4258;
wire net_8371;
wire net_7443;
wire net_12838;
wire net_12454;
wire net_9985;
wire net_13833;
wire net_7301;
wire net_1555;
wire net_10594;
wire net_9349;
wire net_4480;
wire net_10131;
wire net_15454;
wire net_15153;
wire net_2171;
wire net_10233;
wire net_6338;
wire net_18025;
wire net_4521;
wire net_6112;
wire net_2425;
wire net_11245;
wire net_13691;
wire net_18209;
wire net_8319;
wire x3685;
wire net_10573;
wire net_2509;
wire x13534;
wire net_17075;
wire net_2156;
wire net_9177;
wire net_14188;
wire net_8488;
wire net_6831;
wire net_13246;
wire net_4314;
wire net_11640;
wire net_10005;
wire net_3343;
wire net_18188;
wire net_3326;
wire net_11877;
wire net_2239;
wire net_16838;
wire net_3394;
wire net_12846;
wire net_17026;
wire net_4680;
wire net_18595;
wire net_3903;
wire net_15192;
wire net_8879;
wire net_4050;
wire net_16818;
wire net_1571;
wire net_11467;
wire net_16155;
wire net_9248;
wire net_18887;
wire net_5090;
wire net_10530;
wire net_850;
wire net_12511;
wire net_1168;
wire net_10118;
wire net_11008;
wire net_5545;
wire net_9631;
wire net_17685;
wire net_10744;
wire net_3090;
wire net_8747;
wire net_15052;
wire net_8387;
wire net_1009;
wire net_715;
wire net_11444;
wire net_18502;
wire net_13857;
wire net_14503;
wire net_16475;
wire net_8454;
wire net_16152;
wire net_2546;
wire net_11181;
wire net_7056;
wire net_12042;
wire net_15876;
wire net_16810;
wire net_6702;
wire net_312;
wire net_11130;
wire net_2627;
wire net_5386;
wire net_147;
wire net_17237;
wire net_7182;
wire net_12490;
wire net_16453;
wire net_8589;
wire net_12137;
wire x1575;
wire net_7750;
wire net_12335;
wire net_2444;
wire net_17454;
wire net_13496;
wire net_5297;
wire net_8148;
wire net_12936;
wire net_9625;
wire net_17753;
wire net_10122;
wire net_14965;
wire net_8551;
wire net_10759;
wire net_14148;
wire x871;
wire net_7431;
wire net_5398;
wire net_18200;
wire net_2435;
wire net_245;
wire net_6990;
wire net_4858;
wire net_2383;
wire net_12177;
wire net_3491;
wire net_11013;
wire net_16296;
wire net_10829;
wire net_8380;
wire net_277;
wire net_16795;
wire net_4251;
wire net_1965;
wire net_13886;
wire net_680;
wire net_16537;
wire net_17585;
wire net_338;
wire net_13230;
wire net_13435;
wire net_4494;
wire net_8397;
wire net_15672;
wire net_14597;
wire net_9971;
wire net_4089;
wire net_10705;
wire net_13721;
wire net_2009;
wire net_18134;
wire net_17604;
wire net_4026;
wire net_6697;
wire net_1380;
wire net_14844;
wire net_14731;
wire net_9340;
wire net_5176;
wire net_5936;
wire net_18890;
wire net_11956;
wire net_8937;
wire net_6987;
wire net_18469;
wire net_14550;
wire net_1997;
wire net_13206;
wire net_14657;
wire net_15931;
wire net_7718;
wire net_8553;
wire net_6728;
wire net_13364;
wire net_13698;
wire net_11139;
wire net_18897;
wire net_14151;
wire net_6579;
wire net_15232;
wire net_14792;
wire net_1418;
wire net_8686;
wire net_13955;
wire net_5938;
wire net_6980;
wire net_5931;
wire net_8343;
wire net_15226;
wire net_1713;
wire net_12913;
wire net_4684;
wire net_11383;
wire net_8988;
wire net_2775;
wire net_7001;
wire net_14594;
wire net_12007;
wire net_17919;
wire net_14839;
wire net_7654;
wire net_163;
wire net_6022;
wire x13826;
wire net_5802;
wire net_15736;
wire net_11037;
wire net_8037;
wire net_15843;
wire net_19046;
wire net_8444;
wire net_9830;
wire net_18169;
wire net_6135;
wire net_11580;
wire net_13863;
wire net_2193;
wire net_12595;
wire net_12002;
wire net_12293;
wire net_11159;
wire net_18102;
wire net_6304;
wire net_5574;
wire net_11704;
wire net_5258;
wire net_17133;
wire net_1886;
wire x13364;
wire net_2604;
wire net_13689;
wire net_12191;
wire net_14115;
wire net_4678;
wire net_18593;
wire net_14307;
wire net_14256;
wire net_4866;
wire net_5652;
wire net_16256;
wire net_2109;
wire net_1770;
wire net_9326;
wire net_4703;
wire net_17302;
wire net_14530;
wire x13560;
wire net_4770;
wire net_7770;
wire net_378;
wire net_14049;
wire net_14262;
wire net_3309;
wire net_5767;
wire net_16972;
wire net_10032;
wire net_18377;
wire net_4202;
wire net_11628;
wire net_18535;
wire net_1958;
wire net_1931;
wire net_15493;
wire net_14041;
wire net_1549;
wire net_6244;
wire net_10039;
wire net_16883;
wire net_7736;
wire net_2929;
wire net_7192;
wire net_16608;
wire net_7213;
wire net_5666;
wire net_8527;
wire net_11227;
wire net_818;
wire net_15103;
wire net_11275;
wire net_16855;
wire net_1211;
wire net_5448;
wire net_1183;
wire net_4248;
wire net_14537;
wire net_12337;
wire net_17979;
wire net_7241;
wire net_16035;
wire net_17190;
wire net_9753;
wire net_4674;
wire net_9203;
wire net_9551;
wire net_15495;
wire net_6791;
wire net_2017;
wire net_5154;
wire net_11508;
wire net_16138;
wire net_2735;
wire net_12145;
wire net_8780;
wire net_8377;
wire net_16466;
wire net_8800;
wire net_18747;
wire net_1621;
wire net_14432;
wire net_16661;
wire net_18247;
wire net_1035;
wire net_12253;
wire net_11331;
wire net_14076;
wire net_17509;
wire net_13035;
wire net_5597;
wire net_6914;
wire net_4656;
wire net_3593;
wire net_10264;
wire net_6748;
wire net_2641;
wire net_16584;
wire net_7711;
wire net_18972;
wire net_6688;
wire net_9389;
wire net_4035;
wire net_12321;
wire net_18058;
wire net_7816;
wire net_9362;
wire net_9881;
wire net_17697;
wire net_8948;
wire net_9092;
wire net_13464;
wire net_7919;
wire net_2882;
wire net_8131;
wire net_14440;
wire net_14191;
wire net_18785;
wire net_14253;
wire net_3064;
wire net_5731;
wire net_2276;
wire net_6369;
wire net_12748;
wire net_9302;
wire net_11639;
wire net_7748;
wire net_9426;
wire net_6745;
wire net_13716;
wire net_798;
wire net_14149;
wire net_14820;
wire net_18612;
wire net_2059;
wire net_16002;
wire net_18911;
wire net_15806;
wire net_15993;
wire net_9740;
wire net_8520;
wire net_6018;
wire net_8860;
wire net_1336;
wire net_16074;
wire net_18905;
wire net_9915;
wire net_10033;
wire net_6946;
wire x4455;
wire net_11739;
wire net_14114;
wire net_11534;
wire x3996;
wire net_11671;
wire net_3336;
wire net_903;
wire net_9561;
wire net_15502;
wire net_10025;
wire net_12069;
wire net_13796;
wire net_7354;
wire net_8407;
wire net_11395;
wire net_18387;
wire net_5986;
wire net_2378;
wire net_16896;
wire net_17290;
wire net_6261;
wire net_10461;
wire net_11758;
wire net_10319;
wire net_8046;
wire net_17974;
wire net_18238;
wire net_13746;
wire net_15378;
wire net_7125;
wire net_16393;
wire net_8605;
wire net_9865;
wire net_10010;
wire net_14445;
wire net_5566;
wire net_5281;
wire net_8776;
wire net_2327;
wire net_1003;
wire net_8772;
wire net_10868;
wire net_17559;
wire net_15443;
wire net_17552;
wire net_7376;
wire net_11255;
wire net_10310;
wire net_14093;
wire net_5669;
wire net_6122;
wire net_6497;
wire net_6060;
wire net_11991;
wire net_13387;
wire net_16287;
wire net_11513;
wire net_13554;
wire net_3742;
wire net_445;
wire net_13398;
wire net_10773;
wire net_6673;
wire net_12319;
wire net_13637;
wire net_17828;
wire net_18583;
wire net_2213;
wire net_8307;
wire net_2575;
wire net_11986;
wire net_15880;
wire net_9219;
wire net_19006;
wire net_12142;
wire net_6921;
wire net_17099;
wire net_8445;
wire net_13517;
wire net_3713;
wire net_10876;
wire net_556;
wire net_18311;
wire net_4121;
wire x2746;
wire net_3826;
wire net_620;
wire net_18157;
wire net_8702;
wire net_16096;
wire net_4659;
wire net_7321;
wire net_14529;
wire net_5997;
wire net_4779;
wire net_14392;
wire net_16954;
wire net_11150;
wire net_8156;
wire net_5129;
wire net_10444;
wire net_7883;
wire net_17471;
wire net_6414;
wire net_5393;
wire net_17327;
wire net_6937;
wire net_7825;
wire net_13613;
wire net_8855;
wire net_1493;
wire net_17407;
wire x3327;
wire net_9167;
wire net_17459;
wire net_11143;
wire net_8498;
wire net_8897;
wire net_4179;
wire net_2579;
wire net_8235;
wire net_9581;
wire net_6013;
wire net_10296;
wire net_7307;
wire net_5873;
wire net_1866;
wire net_12990;
wire net_14852;
wire net_6934;
wire net_5761;
wire net_3211;
wire net_16552;
wire net_10820;
wire net_13060;
wire net_16798;
wire net_7634;
wire net_5927;
wire net_13894;
wire net_11738;
wire net_12754;
wire net_8625;
wire net_16680;
wire net_8342;
wire net_11732;
wire net_2516;
wire net_18480;
wire net_7553;
wire net_2807;
wire net_4687;
wire net_10676;
wire net_15908;
wire net_18694;
wire net_16655;
wire net_18342;
wire net_6321;
wire net_7584;
wire net_1288;
wire net_16382;
wire net_4708;
wire net_10511;
wire net_12554;
wire net_10559;
wire net_2300;
wire net_8119;
wire net_6710;
wire net_8426;
wire net_7091;
wire net_6383;
wire net_13915;
wire net_6434;
wire net_4816;
wire x364;
wire net_11428;
wire net_11604;
wire net_17760;
wire net_17058;
wire net_5524;
wire net_16381;
wire net_4937;
wire net_4199;
wire net_1043;
wire net_11897;
wire net_16543;
wire net_15086;
wire net_18764;
wire net_18846;
wire net_9737;
wire net_6389;
wire net_16806;
wire net_7493;
wire net_1630;
wire x12922;
wire net_2956;
wire net_18094;
wire net_1082;
wire net_11170;
wire net_15645;
wire net_10405;
wire net_16516;
wire net_16365;
wire net_15407;
wire net_18282;
wire net_11861;
wire net_3296;
wire net_257;
wire net_8543;
wire net_10096;
wire net_11407;
wire net_5500;
wire net_9978;
wire net_5770;
wire net_18682;
wire net_6576;
wire net_958;
wire net_12646;
wire net_4556;
wire net_6400;
wire net_11447;
wire net_12407;
wire net_6199;
wire net_1734;
wire net_10189;
wire net_17205;
wire net_11175;
wire net_5534;
wire net_4308;
wire net_10987;
wire net_17927;
wire net_17041;
wire net_16424;
wire net_7166;
wire net_13450;
wire net_14510;
wire net_3050;
wire net_1728;
wire net_5963;
wire net_12883;
wire net_15394;
wire net_3956;
wire net_16441;
wire net_12426;
wire net_10218;
wire net_8467;
wire net_8761;
wire net_425;
wire net_17818;
wire net_5204;
wire net_17417;
wire net_2205;
wire net_13154;
wire net_8108;
wire net_16123;
wire net_11344;
wire net_17621;
wire net_13667;
wire net_16087;
wire net_368;
wire net_8064;
wire net_4833;
wire net_15914;
wire net_10670;
wire net_2000;
wire net_13089;
wire net_6226;
wire net_14799;
wire net_12502;
wire net_18313;
wire net_2984;
wire net_1020;
wire net_10603;
wire net_15971;
wire net_18366;
wire net_3282;
wire net_3122;
wire net_13989;
wire net_17860;
wire net_8546;
wire net_10164;
wire net_10763;
wire net_16990;
wire net_8594;
wire net_12521;
wire net_18562;
wire net_2094;
wire net_11965;
wire net_7282;
wire net_2543;
wire net_8275;
wire net_760;
wire net_2083;
wire net_8318;
wire net_12050;
wire net_17223;
wire net_3851;
wire net_2488;
wire net_4536;
wire net_5034;
wire net_8192;
wire net_17767;
wire net_1870;
wire net_5200;
wire net_12772;
wire net_2063;
wire net_192;
wire net_17922;
wire net_1739;
wire net_2912;
wire net_4140;
wire net_18293;
wire x1467;
wire net_13254;
wire net_735;
wire net_14269;
wire net_17060;
wire net_3809;
wire net_16824;
wire net_9442;
wire net_1081;
wire net_17636;
wire net_2037;
wire net_8163;
wire net_1237;
wire net_1420;
wire net_12478;
wire net_4789;
wire net_9112;
wire net_14921;
wire net_4064;
wire net_9587;
wire net_4237;
wire net_9712;
wire net_9542;
wire net_17486;
wire net_4559;
wire net_18265;
wire net_7782;
wire net_3144;
wire net_699;
wire net_359;
wire net_5239;
wire net_16940;
wire net_16065;
wire net_9068;
wire net_12862;
wire net_5827;
wire net_2819;
wire net_11316;
wire net_15901;
wire net_882;
wire net_15614;
wire net_6433;
wire net_1827;
wire net_14867;
wire net_4109;
wire net_12606;
wire net_15958;
wire net_8903;
wire net_3858;
wire net_7838;
wire net_10813;
wire net_14182;
wire net_16626;
wire net_15254;
wire net_2283;
wire net_1207;
wire net_10436;
wire net_2121;
wire net_8228;
wire net_14326;
wire net_14671;
wire net_2252;
wire net_4755;
wire net_18733;
wire net_7951;
wire net_17394;
wire net_2126;
wire net_5022;
wire net_9931;
wire net_10449;
wire net_7342;
wire net_16947;
wire net_17657;
wire net_9524;
wire net_12461;
wire net_17398;
wire net_14616;
wire net_18944;
wire net_6952;
wire net_3655;
wire net_17432;
wire net_2304;
wire net_14098;
wire net_12942;
wire net_7418;
wire net_1593;
wire net_8918;
wire net_3380;
wire x12929;
wire net_10397;
wire net_16177;
wire net_15272;
wire net_18511;
wire net_12794;
wire x2908;
wire net_14758;
wire net_11762;
wire x4771;
wire net_5115;
wire net_14682;
wire net_4502;
wire x480;
wire net_15658;
wire net_16844;
wire net_12275;
wire net_2076;
wire net_12567;
wire net_13131;
wire net_6505;
wire net_4378;
wire net_2218;
wire net_6807;
wire net_10147;
wire net_15219;
wire net_1078;
wire net_9811;
wire net_12340;
wire net_9853;
wire net_6813;
wire net_14984;
wire net_6382;
wire net_14896;
wire net_5681;
wire net_13126;
wire x13586;
wire net_10635;
wire net_18930;
wire net_14341;
wire net_12269;
wire net_5197;
wire net_12703;
wire net_13059;
wire net_2355;
wire net_12856;
wire net_13825;
wire net_3262;
wire net_4495;
wire net_12587;
wire net_16438;
wire net_12824;
wire net_7454;
wire net_16379;
wire net_4196;
wire net_3974;
wire net_13678;
wire net_4626;
wire x3891;
wire net_8532;
wire net_8478;
wire net_2976;
wire net_15007;
wire net_13138;
wire net_988;
wire net_8221;
wire net_3621;
wire net_9820;
wire net_12441;
wire net_18917;
wire net_4091;
wire net_17448;
wire net_12110;
wire net_18714;
wire net_2838;
wire net_5614;
wire net_5219;
wire net_1841;
wire net_1249;
wire net_17799;
wire net_4601;
wire net_18791;
wire net_7973;
wire net_3163;
wire net_4928;
wire net_18479;
wire net_6221;
wire net_4417;
wire net_7145;
wire net_822;
wire net_7084;
wire net_15369;
wire net_15523;
wire net_17985;
wire x521;
wire net_6561;
wire net_16749;
wire net_13470;
wire net_6842;
wire net_15691;
wire net_7701;
wire net_1974;
wire net_8010;
wire net_4963;
wire net_9996;
wire net_11480;
wire net_9021;
wire net_1544;
wire net_15798;
wire net_7366;
wire net_4400;
wire net_10044;
wire net_18362;
wire net_15572;
wire net_10340;
wire net_17645;
wire net_7929;
wire net_1174;
wire net_15168;
wire net_6731;
wire net_6664;
wire net_1109;
wire net_12326;
wire net_4224;
wire net_13733;
wire net_3457;
wire net_9683;
wire net_10963;
wire net_5276;
wire net_11721;
wire net_4471;
wire net_1102;
wire net_16861;
wire net_5487;
wire net_13644;
wire net_4976;
wire net_5640;
wire net_5245;
wire net_18928;
wire net_18002;
wire net_11205;
wire net_18622;
wire net_14175;
wire net_2692;
wire net_3777;
wire net_11322;
wire net_18144;
wire net_14355;
wire net_13353;
wire net_10285;
wire net_6279;
wire net_14382;
wire net_15934;
wire net_7516;
wire net_7037;
wire net_1487;
wire net_4572;
wire net_2759;
wire net_10020;
wire net_5408;
wire net_8243;
wire net_3634;
wire net_12486;
wire net_14128;
wire net_13348;
wire net_16570;
wire net_16117;
wire net_18533;
wire net_13705;
wire net_14215;
wire net_10338;
wire net_18650;
wire net_10349;
wire net_2564;
wire net_2821;
wire net_1658;
wire net_5688;
wire net_5481;
wire net_17891;
wire net_7318;
wire net_17823;
wire net_3007;
wire net_7554;
wire net_9505;
wire net_4487;
wire net_15412;
wire net_14998;
wire net_3174;
wire net_9122;
wire net_6966;
wire net_2876;
wire net_844;
wire net_1496;
wire net_325;
wire net_14470;
wire net_1820;
wire net_8175;
wire net_14628;
wire net_5690;
wire net_13274;
wire net_10287;
wire net_16783;
wire net_5956;
wire net_5014;
wire net_7517;
wire net_4036;
wire net_11266;
wire net_1521;
wire net_6274;
wire net_4182;
wire x626;
wire net_11813;
wire net_7908;
wire net_11727;
wire net_7179;
wire net_4734;
wire net_2991;
wire net_4276;
wire net_564;
wire net_10077;
wire net_14919;
wire net_6154;
wire net_10618;
wire net_2050;
wire net_4086;
wire net_9082;
wire net_13992;
wire net_813;
wire net_14105;
wire net_5609;
wire net_10661;
wire net_15279;
wire net_1027;
wire net_1408;
wire net_12403;
wire net_265;
wire net_15819;
wire net_8110;
wire net_11720;
wire net_8673;
wire net_11097;
wire net_13538;
wire net_6774;
wire net_10834;
wire net_9351;
wire net_1155;
wire net_9258;
wire net_14606;
wire net_9787;
wire net_7374;
wire net_12764;
wire net_16324;
wire net_864;
wire net_10331;
wire net_17186;
wire net_7691;
wire net_18569;
wire net_16340;
wire net_13004;
wire net_12787;
wire net_12285;
wire net_16706;
wire net_4113;
wire net_14992;
wire net_17148;
wire net_8850;
wire net_10365;
wire net_16591;
wire net_2298;
wire net_660;
wire net_14060;
wire net_9707;
wire net_6580;
wire net_1908;
wire net_7647;
wire net_9309;
wire net_3383;
wire net_18552;
wire net_13020;
wire net_7265;
wire net_12958;
wire net_6751;
wire net_3914;
wire net_7607;
wire net_6531;
wire net_17084;
wire net_14104;
wire net_6463;
wire net_11973;
wire net_6455;
wire net_5777;
wire net_10610;
wire net_7576;
wire net_13449;
wire net_16595;
wire net_16916;
wire net_2145;
wire net_6488;
wire net_16529;
wire net_11109;
wire net_17101;
wire net_3311;
wire net_8874;
wire net_11020;
wire net_12729;
wire net_14036;
wire net_10887;
wire net_10454;
wire net_15310;
wire net_10716;
wire net_18346;
wire net_4853;
wire net_13943;
wire net_8699;
wire net_14775;
wire net_10474;
wire net_13080;
wire net_3538;
wire net_11507;
wire net_17200;
wire net_17617;
wire net_1583;
wire net_15564;
wire net_9454;
wire net_4408;
wire net_1563;
wire net_3898;
wire net_4948;
wire net_13969;
wire net_7600;
wire net_16349;
wire net_5599;
wire net_13073;
wire net_3361;
wire net_10553;
wire net_13019;
wire net_8578;
wire net_14285;
wire net_15892;
wire net_18255;
wire net_1942;
wire net_11484;
wire net_10070;
wire net_12119;
wire net_13755;
wire net_7891;
wire net_18601;
wire net_1267;
wire net_14150;
wire net_6093;
wire net_3944;
wire net_3661;
wire net_11846;
wire net_12570;
wire net_9188;
wire net_4893;
wire net_18221;
wire net_12982;
wire net_6526;
wire net_5888;
wire net_5131;
wire net_2349;
wire net_18868;
wire net_11074;
wire net_1294;
wire net_10350;
wire net_14450;
wire net_14692;
wire net_3520;
wire net_5006;
wire net_18877;
wire net_1354;
wire net_15480;
wire net_2904;
wire net_1308;
wire net_7631;
wire net_18426;
wire net_4332;
wire net_12081;
wire net_15998;
wire net_1389;
wire net_9992;
wire net_12114;
wire net_13818;
wire net_4748;
wire net_3250;
wire net_5304;
wire net_10737;
wire net_17723;
wire net_548;
wire net_16931;
wire net_4985;
wire net_2402;
wire net_6529;
wire net_5902;
wire net_5082;
wire net_636;
wire net_10239;
wire net_4269;
wire net_18803;
wire net_8159;
wire net_18494;
wire net_8218;
wire net_8471;
wire net_17947;
wire net_12678;
wire net_4262;
wire net_4165;
wire net_16230;
wire net_4506;
wire net_1185;
wire net_10228;
wire net_13868;
wire net_5001;
wire x3258;
wire net_16881;
wire net_7942;
wire net_11216;
wire net_9401;
wire net_4826;
wire net_1912;
wire net_9566;
wire net_11263;
wire net_11353;
wire net_17092;
wire net_11416;
wire net_9118;
wire net_11542;
wire net_9906;
wire net_15746;
wire net_15721;
wire net_18670;
wire net_1538;
wire net_14228;
wire net_9501;
wire net_11499;
wire net_13965;
wire net_1579;
wire net_13440;
wire net_6484;
wire net_10520;
wire net_1999;
wire net_6669;
wire net_1014;
wire net_1444;
wire net_2679;
wire net_17450;
wire net_6255;
wire net_4082;
wire net_11577;
wire net_14666;
wire net_538;
wire net_9083;
wire net_14746;
wire net_14864;
wire net_4130;
wire net_12994;
wire net_9965;
wire net_13306;
wire net_366;
wire net_1854;
wire net_1917;
wire net_1755;
wire net_1359;
wire net_16113;
wire net_2460;
wire net_8929;
wire net_13228;
wire net_14704;
wire net_11238;
wire net_15547;
wire net_11348;
wire net_13424;
wire net_12618;
wire net_14496;
wire net_209;
wire net_1282;
wire net_9242;
wire net_17804;
wire net_17883;
wire net_8211;
wire net_4041;
wire net_13291;
wire net_3204;
wire net_16406;
wire net_8996;
wire net_12315;
wire net_3471;
wire net_18723;
wire net_9677;
wire net_9692;
wire net_12354;
wire net_12966;
wire net_3512;
wire net_15387;
wire x13815;
wire net_8907;
wire net_9394;
wire net_11531;
wire net_10382;
wire net_2430;
wire x406;
wire net_10177;
wire net_4461;
wire net_8433;
wire net_17267;
wire net_7687;
wire net_13598;
wire net_3481;
wire net_11942;
wire net_1589;
wire net_14979;
wire net_17543;
wire net_8114;
wire net_2396;
wire net_9098;
wire net_19032;
wire net_13298;
wire net_15489;
wire net_16771;
wire net_8354;
wire net_5815;
wire net_2856;
wire net_787;
wire net_7777;
wire net_10789;
wire net_8125;
wire net_3603;
wire net_9656;
wire net_16029;
wire net_4187;
wire net_8095;
wire net_16491;
wire net_12071;
wire net_14323;
wire net_8463;
wire net_11001;
wire net_6195;
wire net_10767;
wire net_3579;
wire net_16146;
wire net_18575;
wire net_11069;
wire net_8870;
wire net_2139;
wire net_15638;
wire net_5332;
wire net_10250;
wire net_18633;
wire net_1910;
wire net_8103;
wire net_17158;
wire net_12689;
wire net_14891;
wire net_3544;
wire net_5229;
wire net_3034;
wire net_9517;
wire x12843;
wire net_7895;
wire net_9488;
wire net_7938;
wire net_7610;
wire net_6285;
wire net_18866;
wire net_12817;
wire net_11030;
wire net_2493;
wire net_9664;
wire net_919;
wire net_11914;
wire net_9009;
wire net_11574;
wire net_7044;
wire net_6836;
wire net_6444;
wire net_4008;
wire net_12669;
wire net_15280;
wire net_2209;
wire net_1372;
wire net_1757;
wire net_11935;
wire net_15601;
wire net_5215;
wire net_8816;
wire net_13084;
wire net_13015;
wire net_14547;
wire net_2682;
wire net_7151;
wire net_14936;
wire net_8053;
wire net_17500;
wire net_14562;
wire net_11949;
wire net_6612;
wire net_7077;
wire net_8911;
wire net_3790;
wire net_17313;
wire net_9141;
wire net_15235;
wire net_4267;
wire net_15275;
wire net_12482;
wire net_18394;
wire net_7328;
wire net_2178;
wire net_5292;
wire net_3073;
wire net_10134;
wire net_8840;
wire net_7949;
wire net_13846;
wire net_18420;
wire net_804;
wire net_10541;
wire net_3548;
wire net_1314;
wire net_9400;
wire net_6325;
wire net_8845;
wire net_5376;
wire net_16484;
wire net_531;
wire net_8582;
wire net_499;
wire net_2752;
wire net_9126;
wire net_10701;
wire net_16165;
wire net_17792;
wire net_9476;
wire net_9699;
wire net_4390;
wire net_3534;
wire net_8027;
wire net_13413;
wire net_17844;
wire net_1765;
wire net_12155;
wire net_8965;
wire net_18290;
wire net_10424;
wire net_14878;
wire net_11231;
wire net_6208;
wire net_6068;
wire net_2774;
wire net_2420;
wire net_12437;
wire net_13410;
wire net_1979;
wire net_5135;
wire net_13927;
wire net_1460;
wire net_1451;
wire net_13978;
wire net_12246;
wire net_18195;
wire net_17460;
wire net_5065;
wire net_5008;
wire net_6619;
wire net_8419;
wire net_15860;
wire net_4803;
wire net_14667;
wire net_17777;
wire net_15682;
wire net_203;
wire net_16890;
wire net_6597;
wire net_14589;
wire net_11071;
wire net_1602;
wire net_12213;
wire net_237;
wire net_613;
wire net_9919;
wire net_13239;
wire net_17561;
wire net_14236;
wire net_1095;
wire net_16070;
wire net_4729;
wire net_578;
wire net_12236;
wire net_15467;
wire net_15460;
wire net_14787;
wire net_16616;
wire net_11288;
wire net_8514;
wire net_18457;
wire net_18053;
wire net_14881;
wire net_2743;
wire net_2159;
wire net_388;
wire net_3647;
wire net_14360;
wire net_536;
wire net_1332;
wire net_17786;
wire net_18458;
wire net_3276;
wire net_10589;
wire net_393;
wire net_11980;
wire net_7468;
wire net_13525;
wire net_9130;
wire net_408;
wire net_10904;
wire net_16101;
wire net_15207;
wire net_16449;
wire net_3246;
wire net_10582;
wire net_1845;
wire net_18543;
wire net_10633;
wire net_12225;
wire net_17273;
wire net_17297;
wire net_9939;
wire net_15969;
wire net_15438;
wire net_3390;
wire net_18740;
wire net_15446;
wire net_2372;
wire net_12579;
wire net_12870;
wire net_868;
wire net_11223;
wire net_10979;
wire net_6079;
wire net_6821;
wire net_13750;
wire net_5029;
wire net_13871;
wire net_270;
wire net_522;
wire net_922;
wire net_2638;
wire net_17318;
wire net_9747;
wire net_13355;
wire net_5429;
wire net_15776;
wire net_4992;
wire net_6140;
wire net_5757;
wire net_2264;
wire net_977;
wire net_11632;
wire net_4780;
wire net_643;
wire net_11278;
wire net_6876;
wire net_6175;
wire net_11165;
wire net_13564;
wire net_15340;
wire net_3587;
wire net_3762;
wire net_10580;
wire net_17348;
wire net_3687;
wire net_10056;
wire net_5307;
wire net_10483;
wire net_12015;
wire net_4920;
wire net_3874;
wire net_2045;
wire net_9357;
wire net_11790;
wire net_11829;
wire net_2869;
wire net_3332;
wire net_3446;
wire net_1892;
wire net_18870;
wire net_1798;
wire net_4427;
wire net_7401;
wire net_13109;
wire net_837;
wire net_13287;
wire net_3469;
wire net_10723;
wire net_9449;
wire net_927;
wire net_11686;
wire net_15838;
wire net_17375;
wire net_693;
wire net_1519;
wire net_12633;
wire net_17992;
wire net_16665;
wire net_6378;
wire net_11390;
wire net_17736;
wire net_3964;
wire net_13777;
wire net_12660;
wire net_4219;
wire net_9311;
wire net_15166;
wire net_9898;
wire net_11865;
wire net_15816;
wire net_14632;
wire net_10847;
wire net_17847;
wire net_13391;
wire net_10208;
wire net_11651;
wire net_488;
wire net_4909;
wire net_10460;
wire net_12009;
wire net_6034;
wire net_18287;
wire net_17170;
wire net_5452;
wire net_8088;
wire net_2319;
wire net_8324;
wire net_15717;
wire net_7102;
wire net_5458;
wire net_11785;
wire net_1532;
wire net_8440;
wire net_8971;
wire net_6653;
wire net_12308;
wire net_4475;
wire net_8207;
wire net_16981;
wire net_11595;
wire net_15478;
wire net_7765;
wire net_14639;
wire net_4958;
wire net_15215;
wire net_14719;
wire net_5057;
wire net_1093;
wire net_2592;
wire net_14947;
wire net_7680;
wire net_6230;
wire net_16343;
wire net_3580;
wire net_9876;
wire net_15505;
wire net_16641;
wire net_3259;
wire net_5260;
wire net_9877;
wire net_10057;
wire net_8833;
wire net_710;
wire net_8922;
wire net_14908;
wire net_17301;
wire net_18020;
wire net_17608;
wire net_14754;
wire net_15072;
wire net_3097;
wire net_14686;
wire net_5836;
wire net_6478;
wire net_16866;
wire net_14401;
wire net_17745;
wire net_18320;
wire net_3970;
wire net_3018;
wire net_173;
wire net_12516;
wire net_14317;
wire net_9237;
wire net_16264;
wire net_6203;
wire net_3006;
wire x13594;
wire net_16778;
wire net_16273;
wire net_10970;
wire net_1681;
wire net_16131;
wire net_7936;
wire net_17632;
wire net_14468;
wire net_7998;
wire net_15511;
wire net_4272;
wire net_16726;
wire net_6512;
wire net_10532;
wire net_746;
wire net_13406;
wire net_6147;
wire net_5877;
wire net_17153;
wire net_1274;
wire net_1682;
wire net_11302;
wire net_5743;
wire net_10788;
wire net_7910;
wire net_14485;
wire net_18555;
wire net_10109;
wire net_3466;
wire net_16623;
wire net_15784;
wire net_4995;
wire net_7834;
wire net_629;
wire net_1663;
wire net_14579;
wire net_4209;
wire net_8666;
wire net_15326;
wire net_9382;
wire net_3019;
wire net_13784;
wire net_15017;
wire net_5579;
wire net_14710;
wire net_2351;
wire net_18950;
wire net_17244;
wire x2355;
wire net_1350;
wire net_9628;
wire net_14457;
wire net_1648;
wire net_6219;
wire net_12594;
wire net_631;
wire net_14201;
wire net_12128;
wire net_16603;
wire net_10086;
wire net_17811;
wire net_14988;
wire net_13143;
wire net_4007;
wire net_4499;
wire net_8566;
wire net_12100;
wire net_9910;
wire net_15733;
wire net_16306;
wire net_6928;
wire net_670;
wire net_15159;
wire net_6250;
wire net_2687;
wire net_9889;
wire net_7023;
wire net_10750;
wire net_9721;
wire net_9842;
wire net_12853;
wire net_16687;
wire net_3928;
wire net_13369;
wire net_14540;
wire net_7038;
wire net_3854;
wire net_6717;
wire net_9793;
wire net_9857;
wire net_5493;
wire net_13759;
wire net_755;
wire net_17522;
wire net_9557;
wire net_7754;
wire net_9285;
wire net_14981;
wire net_12545;
wire net_5892;
wire net_16187;
wire net_13468;
wire net_3151;
wire net_14953;
wire net_6763;
wire net_12890;
wire net_6053;
wire net_3628;
wire net_18778;
wire net_12023;
wire net_18223;
wire net_14479;
wire net_12829;
wire net_16303;
wire net_1652;
wire net_11319;
wire net_16213;
wire net_1429;
wire net_11061;
wire net_14223;
wire net_14895;
wire net_7130;
wire net_18851;
wire net_15223;
wire net_2725;
wire net_3613;
wire net_13166;
wire x1062;
wire net_8964;
wire net_4615;
wire net_727;
wire net_11242;
wire net_9804;
wire net_16259;
wire net_12559;
wire net_4955;
wire net_3190;
wire net_16022;
wire net_3757;
wire net_11457;
wire net_15750;
wire net_18836;
wire net_9224;
wire net_12658;
wire net_4445;
wire net_15142;
wire net_11115;
wire net_14247;
wire net_3951;
wire net_14614;
wire net_15054;
wire net_11635;
wire net_13010;
wire net_2259;
wire net_12124;
wire net_15079;
wire net_10651;
wire net_15107;
wire net_16319;
wire net_4095;
wire net_2739;
wire net_13330;
wire net_10113;
wire net_11715;
wire net_2110;
wire net_2919;
wire net_10642;
wire net_2893;
wire net_11435;
wire net_3227;
wire net_2358;
wire net_16335;
wire net_17465;
wire net_12651;
wire net_8682;
wire net_3057;
wire net_9039;
wire net_571;
wire net_10692;
wire net_10543;
wire net_7569;
wire net_16719;
wire net_14743;
wire net_10400;
wire net_4935;
wire net_3934;
wire net_12168;
wire net_17938;
wire net_10385;
wire net_1877;
wire net_720;
wire net_16107;
wire net_7653;
wire net_9038;
wire net_12152;
wire net_15978;
wire net_18752;
wire net_14005;
wire net_18509;
wire net_5209;
wire net_2199;
wire net_10628;
wire net_684;
wire net_2648;
wire net_16414;
wire net_7299;
wire net_7542;
wire net_3720;
wire net_510;
wire net_12922;
wire net_10909;
wire net_15808;
wire x13508;
wire net_8885;
wire net_2653;
wire net_2960;
wire net_9078;
wire net_8257;
wire net_6703;
wire net_12577;
wire net_7043;
wire net_2782;
wire net_494;
wire net_17364;
wire net_17693;
wire net_10999;
wire net_12877;
wire net_4283;
wire net_15726;
wire net_6592;
wire net_13830;
wire net_18095;
wire net_6084;
wire net_8953;
wire net_16044;
wire net_3461;
wire net_12365;
wire net_10327;
wire net_10956;
wire net_11747;
wire net_4610;
wire net_14366;
wire net_4459;
wire net_457;
wire net_2246;
wire net_8821;
wire net_12096;
wire net_772;
wire net_10180;
wire net_4371;
wire net_14375;
wire net_10190;
wire net_12773;
wire net_7966;
wire net_11807;
wire net_1277;
wire net_14567;
wire net_17712;
wire net_2661;
wire net_16496;
wire net_6113;
wire net_3893;
wire net_13459;
wire net_18988;
wire net_12467;
wire net_4075;
wire net_6421;
wire net_7385;
wire net_18589;
wire net_6051;
wire net_2852;
wire net_1721;
wire net_7851;
wire net_16370;
wire net_12975;
wire net_4633;
wire net_6605;
wire net_6249;
wire net_5843;
wire net_10626;
wire net_1073;
wire net_8073;
wire net_18064;
wire net_17626;
wire net_1947;
wire net_11932;
wire net_879;
wire net_7227;
wire net_2415;
wire net_15034;
wire net_8738;
wire net_7312;
wire net_13225;
wire net_3197;
wire net_1348;
wire net_10740;
wire net_15707;
wire net_17371;
wire net_9774;
wire net_7276;
wire net_16997;
wire net_17388;
wire net_7201;
wire net_18781;
wire net_16017;
wire x13633;
wire net_3422;
wire net_199;
wire net_10151;
wire net_2789;
wire net_7844;
wire net_16397;
wire net_3835;
wire net_431;
wire net_12903;
wire net_5783;
wire net_8250;
wire net_17874;
wire net_9373;
wire net_10898;
wire net_5186;
wire net_4362;
wire net_222;
wire net_13215;
wire net_17255;
wire net_4520;
wire net_15727;
wire net_7804;
wire net_7060;
wire net_3999;
wire net_1788;
wire net_16694;
wire net_4301;
wire net_12476;
wire net_2935;
wire net_6166;
wire net_18841;
wire net_4345;
wire net_10507;
wire net_9318;
wire net_3516;
wire net_6547;
wire net_11799;
wire net_4588;
wire net_1438;
wire net_10374;
wire net_4395;
wire net_8502;
wire net_1143;
wire net_14580;
wire net_15884;
wire net_1088;
wire net_6410;
wire net_9434;
wire net_13262;
wire net_3885;
wire net_706;
wire net_18015;
wire net_6373;
wire net_9298;
wire net_14376;
wire net_2768;
wire net_5125;
wire net_17575;
wire net_551;
wire net_12536;
wire net_13479;
wire net_5368;
wire net_7873;
wire net_4617;
wire net_13182;
wire net_15000;
wire net_11033;
wire net_4168;
wire net_12419;
wire x789;
wire net_12376;
wire net_16979;
wire net_1199;
wire net_11371;
wire net_18081;
wire net_7986;
wire net_8930;
wire net_15675;
wire net_3627;
wire net_14764;
wire net_18032;
wire net_15087;
wire net_5530;
wire net_15296;
wire net_4869;
wire net_450;
wire net_289;
wire net_19021;
wire net_8041;
wire net_9046;
wire net_14204;
wire net_10972;
wire net_2614;
wire net_1642;
wire net_12158;
wire net_5322;
wire net_16958;
wire net_2524;
wire net_11490;
wire net_1224;
wire net_6786;
wire net_13804;
wire net_768;
wire net_11084;
wire net_14423;
wire net_14068;
wire net_908;
wire net_19028;
wire net_18969;
wire net_13189;
wire net_519;
wire x13994;
wire net_9697;
wire net_11773;
wire net_11052;
wire net_2697;
wire net_15825;
wire net_9184;
wire net_10808;
wire x13433;
wire net_6282;
wire net_1204;
wire net_9190;
wire net_14082;
wire net_18216;
wire net_16312;
wire net_14089;
wire net_16923;
wire net_2342;
wire net_7336;
wire net_8331;
wire net_6628;
wire net_9969;
wire net_18719;
wire net_6778;
wire net_3214;
wire net_1986;
wire net_16679;
wire net_14972;
wire net_11472;
wire net_10864;
wire net_12881;
wire net_18405;
wire net_15321;
wire net_6467;
wire net_8203;
wire net_16528;
wire net_7527;
wire net_12613;
wire net_3406;
wire net_9012;
wire net_9164;
wire net_11657;
wire net_4229;
wire net_13110;
wire net_15624;
wire net_6474;
wire net_2130;
wire net_3362;
wire net_1148;
wire net_10198;
wire net_2382;
wire net_13620;
wire net_10698;
wire net_3442;
wire net_5942;
wire net_3864;
wire net_9271;
wire net_15357;
wire net_17063;
wire net_5796;
wire net_9730;
wire net_14725;
wire net_9416;
wire net_6975;
wire net_16355;
wire net_4389;
wire net_11798;
wire net_13935;
wire net_10728;
wire net_10425;
wire net_4561;
wire net_11676;
wire net_14800;
wire net_1473;
wire net_15964;
wire net_1674;
wire net_5582;
wire net_1651;
wire net_2375;
wire net_5109;
wire net_13582;
wire net_6422;
wire net_1806;
wire net_3234;
wire net_15666;
wire net_17578;
wire net_17211;
wire net_8746;
wire net_1363;
wire net_1869;
wire net_4053;
wire net_10526;
wire net_13029;
wire net_15713;
wire net_19018;
wire net_16863;
wire net_4012;
wire net_6169;
wire net_18975;
wire net_6647;
wire net_18503;
wire net_3681;
wire net_6621;
wire net_7902;
wire net_13097;
wire net_7503;
wire net_7857;
wire net_12717;
wire net_10015;
wire net_14522;
wire net_15180;
wire net_5246;
wire net_17982;
wire net_351;
wire net_8558;
wire net_7761;
wire net_12601;
wire net_6006;
wire net_10856;
wire net_4240;
wire net_7964;
wire net_15581;
wire net_2842;
wire net_3158;
wire net_1257;
wire net_939;
wire net_8365;
wire net_18810;
wire net_17424;
wire x420;
wire net_13781;
wire net_7984;
wire net_14411;
wire net_2791;
wire net_10479;
wire net_10111;
wire net_16513;
wire net_11023;
wire net_4271;
wire net_8795;
wire net_15047;
wire net_9895;
wire net_11817;
wire net_317;
wire net_856;
wire net_17001;
wire net_11853;
wire net_9944;
wire net_7920;
wire net_3845;
wire net_16756;
wire net_2026;
wire net_16209;
wire net_5727;
wire net_11822;
wire net_18004;
wire net_16611;
wire net_5673;
wire net_12195;
wire net_3033;
wire net_16567;
wire net_14059;
wire net_18931;
wire net_17037;
wire net_3373;
wire net_5382;
wire net_17854;
wire net_2672;
wire net_11471;
wire net_5351;
wire net_588;
wire net_16648;
wire net_2200;
wire net_8641;
wire net_1157;
wire net_7486;
wire net_7785;
wire net_6001;
wire net_9378;
wire net_14198;
wire net_16922;
wire net_6350;
wire net_7993;
wire net_9840;
wire net_10560;
wire net_14270;
wire net_11800;
wire net_17704;
wire net_13604;
wire net_5603;
wire net_17830;
wire net_1065;
wire net_13117;
wire net_15831;
wire net_3795;
wire net_16245;
wire net_13046;
wire net_16450;
wire net_3100;
wire net_15696;
wire net_13375;
wire net_241;
wire net_9353;
wire net_13196;
wire net_12010;
wire net_13515;
wire net_13640;
wire net_13350;
wire net_4597;
wire net_16291;
wire net_599;
wire net_13814;
wire net_4589;
wire net_4844;
wire net_5860;
wire net_3111;
wire net_18437;
wire net_10346;
wire net_11880;
wire net_13543;
wire net_16765;
wire net_9653;
wire net_8692;
wire net_13575;
wire net_8356;
wire net_18445;
wire net_3737;
wire net_18049;
wire net_6103;
wire net_15384;
wire net_18645;
wire net_12260;
wire net_15752;
wire net_15918;
wire net_9686;
wire net_17141;
wire net_2849;
wire net_12671;
wire net_18638;
wire net_10799;
wire net_15641;
wire net_15267;
wire net_12693;
wire net_5589;
wire net_17535;
wire net_4873;
wire net_10851;
wire net_16461;
wire net_4298;
wire net_16564;
wire net_11286;
wire net_15175;
wire net_18812;
wire net_16876;
wire net_7170;
wire net_8004;
wire net_11250;
wire net_4137;
wire net_8528;
wire net_5162;
wire net_9870;
wire net_17545;
wire net_7561;
wire net_5765;
wire net_3496;
wire net_15010;
wire net_4216;
wire net_13361;
wire net_4889;
wire x1087;
wire net_10371;
wire net_151;
wire net_16950;
wire net_1625;
wire net_13638;
wire net_8784;
wire net_9930;
wire net_17915;
wire net_2513;
wire net_8662;
wire net_7360;
wire net_7142;
wire net_10291;
wire net_187;
wire net_3305;
wire net_14072;
wire net_14045;
wire net_18310;
wire net_160;
wire net_832;
wire net_12304;
wire net_7728;
wire net_6749;
wire net_5578;
wire x4154;
wire net_18659;
wire net_13742;
wire net_6501;
wire net_17868;
wire net_16577;
wire net_9580;
wire net_5272;
wire net_6240;
wire net_7812;
wire net_3838;
wire net_7768;
wire net_11518;
wire net_19031;
wire net_6260;
wire net_15116;
wire net_292;
wire net_12489;
wire net_5529;
wire net_9384;
wire net_12141;
wire net_167;
wire net_12371;
wire net_7308;
wire net_6170;
wire net_8864;
wire net_15325;
wire net_9847;
wire net_15849;
wire net_5735;
wire net_2806;
wire net_9679;
wire net_13163;
wire net_14624;
wire net_4924;
wire net_4483;
wire net_8391;
wire net_9367;
wire net_5045;
wire net_14441;
wire net_17540;
wire net_6237;
wire net_11335;
wire net_2456;
wire net_2753;
wire net_1232;
wire net_10036;
wire net_14635;
wire net_4540;
wire net_9585;
wire net_5662;
wire net_3059;
wire net_11625;
wire net_13506;
wire net_10684;
wire net_12540;
wire net_5444;
wire net_17090;
wire net_13039;
wire net_17436;
wire net_464;
wire net_12003;
wire net_17286;
wire net_5699;
wire net_5089;
wire net_4200;
wire net_6300;
wire net_5867;
wire net_16629;
wire net_5362;
wire net_18539;
wire net_4658;
wire net_12625;
wire net_14195;
wire net_14602;
wire net_1256;
wire net_1413;
wire net_14252;
wire net_15262;
wire net_18997;
wire net_3556;
wire net_1840;
wire net_3041;
wire net_13872;
wire net_12602;
wire net_5637;
wire net_8015;
wire net_7167;
wire net_3427;
wire net_1031;
wire net_13170;
wire net_10265;
wire net_13394;
wire net_7245;
wire net_7458;
wire net_9744;
wire net_10467;
wire net_10991;
wire net_1688;
wire net_2020;
wire net_8523;
wire net_16787;
wire net_15968;
wire net_10794;
wire net_13522;
wire net_7665;
wire net_13383;
wire net_15858;
wire net_6126;
wire net_14056;
wire net_17527;
wire net_15076;
wire net_16684;
wire net_4324;
wire net_4159;
wire net_7322;
wire net_2374;
wire net_4203;
wire net_9911;
wire net_17663;
wire net_10571;
wire net_16039;
wire net_250;
wire net_3600;
wire net_8655;
wire net_7260;
wire net_5882;
wire net_2055;
wire net_12929;
wire net_7420;
wire net_403;
wire net_10027;
wire net_3524;
wire net_6265;
wire net_13680;
wire net_12219;
wire net_15560;
wire net_18699;
wire net_14302;
wire net_9899;
wire net_19000;
wire net_12202;
wire net_12562;
wire net_8602;
wire net_14910;
wire net_794;
wire net_2397;
wire net_8136;
wire net_13277;
wire net_10537;
wire net_3433;
wire net_1468;
wire net_4774;
wire net_11767;
wire net_16360;
wire net_7350;
wire net_8494;
wire net_6796;
wire net_1130;
wire net_5921;
wire net_14826;
wire net_8111;
wire net_8239;
wire net_9421;
wire net_6451;
wire net_7918;
wire net_6493;
wire net_9281;
wire net_7745;
wire net_6309;
wire net_2318;
wire net_8787;
wire net_9207;
wire net_5562;
wire net_17166;
wire net_3449;
wire net_9004;
wire net_9134;
wire net_18463;
wire net_17475;
wire net_1039;
wire net_7822;
wire net_11972;
wire net_4651;
wire net_400;
wire net_8629;
wire net_15499;
wire net_14546;
wire net_1935;
wire net_11608;
wire net_13102;
wire net_2925;
wire net_9142;
wire net_11873;
wire net_18826;
wire net_1855;
wire net_14956;
wire net_4882;
wire net_1163;
wire net_1177;
wire net_10206;
wire net_13890;
wire net_5466;
wire net_9521;
wire net_7840;
wire net_16053;
wire net_17029;
wire net_9215;
wire net_11494;
wire net_3273;
wire net_17978;
wire x933;
wire net_1559;
wire net_5665;
wire net_8706;
wire net_1620;
wire net_2608;
wire net_13966;
wire net_14266;
wire net_2813;
wire net_9763;
wire net_14856;
wire net_14559;
wire net_719;
wire net_10878;
wire net_18234;
wire net_6873;
wire net_8068;
wire net_14032;
wire net_2571;
wire net_9888;
wire net_16892;
wire net_17886;
wire net_16066;
wire net_5703;
wire net_12264;
wire net_9418;
wire net_14325;
wire net_3479;
wire net_8609;
wire net_3222;
wire net_13617;
wire net_16134;
wire net_6393;
wire net_8410;
wire net_3552;
wire net_15314;
wire net_696;
wire net_7427;
wire net_5713;
wire net_10777;
wire net_10824;
wire net_14079;
wire net_17824;
wire net_13175;
wire net_10401;
wire net_13947;
wire net_12972;
wire net_16058;
wire net_12256;
wire net_10448;
wire net_15599;
wire net_9953;
wire net_16093;
wire net_15492;
wire net_17998;
wire net_3821;
wire net_16217;
wire net_9228;
wire net_14101;
wire net_8403;
wire net_4503;
wire net_10872;
wire net_6938;
wire net_3486;
wire net_7359;
wire net_15241;
wire net_17333;
wire net_5839;
wire net_7955;
wire net_8590;
wire net_11199;
wire net_8919;
wire net_9981;
wire net_8302;
wire net_1298;
wire net_296;
wire net_9733;
wire net_16040;
wire net_7004;
wire net_12053;
wire net_18574;
wire net_8941;
wire net_5435;
wire net_17461;
wire net_18071;
wire net_11461;
wire net_18568;
wire net_3020;
wire net_17233;
wire net_13720;
wire net_18205;
wire net_10518;
wire net_1339;
wire net_10608;
wire net_3781;
wire net_17169;
wire net_5685;
wire net_906;
wire net_15450;
wire net_2422;
wire net_5205;
wire net_13951;
wire net_652;
wire net_10185;
wire net_12955;
wire net_13958;
wire net_13707;
wire x13330;
wire net_10590;
wire net_10211;
wire net_14840;
wire net_14513;
wire net_2505;
wire net_11185;
wire net_16988;
wire net_10748;
wire net_6139;
wire net_2683;
wire net_17516;
wire net_4812;
wire net_16180;
wire net_4253;
wire net_2165;
wire net_11943;
wire net_8315;
wire net_6861;
wire net_18821;
wire net_11049;
wire net_2562;
wire net_15417;
wire net_5134;
wire net_5293;
wire net_9129;
wire net_14931;
wire net_7195;
wire net_13841;
wire x1855;
wire net_8151;
wire net_16079;
wire net_5172;
wire net_2182;
wire net_8145;
wire net_10092;
wire net_4718;
wire net_8032;
wire net_9928;
wire net_9295;
wire net_150;
wire net_6589;
wire net_11915;
wire net_16151;
wire net_4351;
wire net_6993;
wire net_10951;
wire net_12436;
wire net_15773;
wire net_7666;
wire net_1703;
wire net_12768;
wire net_11004;
wire net_7848;
wire net_9420;
wire x306;
wire net_9690;
wire net_3693;
wire net_9027;
wire net_5100;
wire net_4319;
wire net_14849;
wire net_18317;
wire net_16246;
wire net_3070;
wire net_13695;
wire net_3409;
wire net_9481;
wire net_17022;
wire net_4525;
wire net_16782;
wire net_1904;
wire net_3907;
wire net_9446;
wire net_6332;
wire net_16493;
wire net_6584;
wire net_10001;
wire net_8617;
wire net_2187;
wire net_17639;
wire net_10764;
wire net_3387;
wire net_13242;
wire net_7157;
wire net_1479;
wire net_16127;
wire net_10268;
wire net_15611;
wire net_18532;
wire net_6895;
wire net_10066;
wire net_3094;
wire net_1927;
wire net_10243;
wire net_213;
wire net_6910;
wire x2041;
wire net_9244;
wire net_947;
wire net_5359;
wire net_7970;
wire net_1126;
wire net_14715;
wire net_2004;
wire net_11538;
wire net_16636;
wire net_6943;
wire net_1325;
wire net_16474;
wire net_5094;
wire net_6298;
wire net_2567;
wire net_10258;
wire net_10944;
wire net_14029;
wire net_7643;
wire net_7411;
wire net_16445;
wire net_1303;
wire net_16158;
wire net_8050;
wire net_18029;
wire net_16834;
wire net_6334;
wire net_18260;
wire net_2102;
wire net_4451;
wire net_1807;
wire net_11903;
wire net_1930;
wire net_1943;
wire net_17493;
wire net_16994;
wire net_17955;
wire net_16471;
wire net_12113;
wire net_4054;
wire net_11555;
wire net_5544;
wire net_18180;
wire net_15842;
wire net_18744;
wire net_5054;
wire net_9674;
wire net_4848;
wire net_7791;
wire net_16114;
wire net_18165;
wire net_3889;
wire net_14899;
wire net_14039;
wire net_3567;
wire net_13717;
wire net_7831;
wire net_11525;
wire net_6483;
wire net_16323;
wire net_6616;
wire net_2448;
wire net_15285;
wire net_5424;
wire net_5541;
wire net_13234;
wire net_10719;
wire net_3400;
wire net_17601;
wire net_14925;
wire net_646;
wire net_5823;
wire net_2731;
wire net_2601;
wire net_11016;
wire net_8902;
wire net_8499;
wire net_520;
wire net_10159;
wire net_13482;
wire net_7237;
wire net_11201;
wire net_4722;
wire net_14110;
wire net_16061;
wire net_3231;
wire net_981;
wire net_18961;
wire net_9636;
wire net_8895;
wire net_1566;
wire net_17941;
wire net_11584;
wire net_2354;
wire net_12156;
wire net_9393;
wire net_10378;
wire net_10709;
wire net_10440;
wire net_5018;
wire net_8858;
wire net_15676;
wire net_7369;
wire net_5013;
wire net_15856;
wire net_559;
wire net_11413;
wire net_16886;
wire net_3042;
wire net_12804;
wire net_7476;
wire net_1717;
wire net_6553;
wire net_398;
wire net_3399;
wire net_6976;
wire net_17072;
wire net_16943;
wire net_6693;
wire net_2117;
wire net_12834;
wire net_4085;
wire net_7393;
wire net_13493;
wire net_10099;
wire net_17797;
wire net_12472;
wire net_18617;
wire net_5905;
wire net_9788;
wire net_15233;
wire net_17589;
wire net_6724;
wire net_6054;
wire net_18845;
wire net_18130;
wire net_1572;
wire net_11647;
wire net_9265;
wire x4570;
wire net_5179;
wire net_2134;
wire net_15595;
wire net_5011;
wire net_316;
wire net_4250;
wire x719;
wire net_13439;
wire net_4961;
wire net_15303;
wire net_4184;
wire net_11462;
wire net_14736;
wire net_14398;
wire net_7033;
wire net_14962;
wire net_17906;
wire net_4647;
wire net_16523;
wire net_4022;
wire net_15649;
wire net_18553;
wire net_17490;
wire net_9618;
wire net_8347;
wire net_13282;
wire net_10040;
wire net_1695;
wire net_5932;
wire net_1617;
wire net_7005;
wire net_5969;
wire net_16815;
wire net_9332;
wire net_18892;
wire net_4579;
wire net_568;
wire net_13809;
wire net_4807;
wire net_1227;
wire net_6046;
wire net_1008;
wire net_5340;
wire net_18848;
wire net_12178;
wire net_4862;
wire net_3069;
wire net_3170;
wire net_12239;
wire x4295;
wire net_4819;
wire net_17613;
wire net_17144;
wire net_14773;
wire net_14533;
wire net_15794;
wire net_469;
wire net_1978;
wire net_18307;
wire net_3167;
wire net_1170;
wire net_5656;
wire net_10144;
wire net_2280;
wire net_13202;
wire net_9174;
wire net_778;
wire net_2366;
wire net_1455;
wire net_2930;
wire net_9816;
wire net_15937;
wire net_14277;
wire net_15651;
wire net_16252;
wire net_16533;
wire net_5323;
wire net_12167;
wire net_6225;
wire net_18654;
wire net_6832;
wire net_5261;
wire net_4730;
wire net_6643;
wire net_11123;
wire net_17505;
wire net_15292;
wire net_4119;
wire net_18148;
wire net_16976;
wire net_9216;
wire net_9450;
wire net_13445;
wire net_18037;
wire net_10335;
wire net_5645;
wire net_995;
wire net_15763;
wire net_8328;
wire net_17790;
wire net_7088;
wire net_7334;
wire net_12232;
wire net_1246;
wire net_8957;
wire net_7705;
wire net_13325;
wire net_1774;
wire net_16162;
wire net_4228;
wire x1174;
wire net_11402;
wire net_3060;
wire net_10712;
wire net_2568;
wire net_11103;
wire net_17008;
wire net_321;
wire net_5518;
wire net_9465;
wire net_17708;
wire net_2995;
wire net_16912;
wire net_3526;
wire net_15532;
wire x778;
wire net_934;
wire net_18795;
wire net_3103;
wire net_5941;
wire net_4896;
wire net_3630;
wire net_11952;
wire net_1824;
wire net_12037;
wire net_7603;
wire net_4763;
wire net_16008;
wire net_5074;
wire net_5694;
wire net_3166;
wire net_18983;
wire net_7065;
wire net_9104;
wire net_8079;
wire net_9831;
wire net_10861;
wire net_7513;
wire net_18272;
wire net_9652;
wire net_10665;
wire net_5552;
wire net_860;
wire net_16566;
wire net_9254;
wire net_2046;
wire net_14474;
wire net_7926;
wire net_11708;
wire net_2878;
wire net_2871;
wire net_9850;
wire net_18325;
wire net_3267;
wire net_2321;
wire net_9108;
wire net_817;
wire net_11667;
wire net_3414;
wire net_15006;
wire net_18349;
wire net_14804;
wire net_7058;
wire net_10967;
wire net_13502;
wire net_9766;
wire net_4576;
wire net_13655;
wire net_13344;
wire net_14123;
wire net_13278;
wire net_5483;
wire net_2012;
wire net_7139;
wire net_5557;
wire net_9890;
wire net_15178;
wire net_16690;
wire net_743;
wire net_3770;
wire net_14387;
wire net_1922;
wire net_9062;
wire net_15333;
wire net_14620;
wire net_17728;
wire net_6639;
wire net_12384;
wire net_8264;
wire net_2451;
wire net_13499;
wire net_14332;
wire net_17012;
wire net_17019;
wire net_4031;
wire net_1522;
wire net_2926;
wire net_12782;
wire net_15881;
wire net_16745;
wire net_8042;
wire net_12289;
wire net_17444;
wire net_13751;
wire net_18883;
wire net_6991;
wire net_4551;
wire net_5972;
wire net_13557;
wire net_18588;
wire net_12945;
wire net_3943;
wire net_9370;
wire net_14996;
wire net_15183;
wire net_17305;
wire net_7675;
wire net_4438;
wire net_10839;
wire net_8557;
wire net_14154;
wire net_968;
wire net_17357;
wire net_13876;
wire net_13572;
wire net_9669;
wire net_10421;
wire net_12692;
wire net_16574;
wire net_17232;
wire net_18416;
wire net_2534;
wire net_6827;
wire net_4133;
wire net_15930;
wire net_3732;
wire net_17835;
wire net_16429;
wire net_2309;
wire net_502;
wire net_8647;
wire net_1564;
wire net_16047;
wire net_6632;
wire net_3804;
wire net_12282;
wire net_10883;
wire net_15353;
wire net_9398;
wire net_17106;
wire net_17046;
wire net_13271;
wire net_8290;
wire net_16707;
wire net_12209;
wire net_13858;
wire net_7990;
wire net_4112;
wire net_3868;
wire net_7121;
wire net_5887;
wire net_13233;
wire net_2628;
wire net_4512;
wire net_6535;
wire net_9305;
wire net_11692;
wire net_17449;
wire net_5145;
wire net_11439;
wire net_12757;
wire net_11160;
wire net_9047;
wire net_10494;
wire net_11078;
wire net_13837;
wire net_13800;
wire net_664;
wire net_6292;
wire net_4622;
wire net_4605;
wire net_4295;
wire net_10450;
wire net_10687;
wire net_12533;
wire net_15684;
wire net_5773;
wire net_10614;
wire net_6405;
wire net_17085;
wire net_18448;
wire net_13550;
wire net_14779;
wire net_7469;
wire net_6210;
wire net_2952;
wire net_2035;
wire net_17429;
wire net_17403;
wire net_5070;
wire net_2826;
wire net_10451;
wire x898;
wire net_17173;
wire net_6847;
wire net_2141;
wire net_15123;
wire net_10830;
wire net_14211;
wire net_11803;
wire net_14818;
wire net_15866;
wire net_19012;
wire net_11213;
wire net_3453;
wire net_5702;
wire net_12648;
wire net_8632;
wire net_9822;
wire net_10598;
wire net_15447;
wire net_6097;
wire net_1403;
wire net_4532;
wire net_2270;
wire net_1667;
wire net_7208;
wire net_8882;
wire net_1606;
wire net_3710;
wire net_15156;
wire net_3054;
wire net_7683;
wire net_17680;
wire net_8765;
wire net_3978;
wire net_16802;
wire net_4752;
wire net_12708;
wire net_15403;
wire net_15704;
wire x4886;
wire net_2029;
wire net_5328;
wire net_3698;
wire net_11560;
wire net_4629;
wire net_2587;
wire net_2959;
wire net_1888;
wire net_11836;
wire net_9974;
wire net_4311;
wire net_18690;
wire net_12583;
wire net_16848;
wire net_1792;
wire net_2496;
wire net_4125;
wire net_17053;
wire net_10656;
wire net_3109;
wire net_1598;
wire net_17390;
wire net_14192;
wire net_731;
wire net_14369;
wire net_17221;
wire net_15063;
wire net_17698;
wire net_15896;
wire net_13042;
wire net_18185;
wire net_7287;
wire net_9704;
wire net_1733;
wire net_5853;
wire net_10576;
wire net_5511;
wire net_7590;
wire net_17737;
wire net_13962;
wire net_11093;
wire net_6708;
wire net_10412;
wire net_18888;
wire net_4146;
wire net_1724;
wire net_6106;
wire net_3703;
wire net_12551;
wire net_17120;
wire net_12682;
wire net_17209;
wire net_12506;
wire net_10843;
wire net_965;
wire net_12378;
wire net_15472;
wire net_17129;
wire net_16457;
wire net_2916;
wire net_5348;
wire net_421;
wire net_8184;
wire net_8314;
wire net_11976;
wire net_1104;
wire net_9783;
wire net_764;
wire net_18120;
wire net_4060;
wire net_5181;
wire net_13009;
wire net_18258;
wire net_5038;
wire net_12465;
wire net_7289;
wire net_1117;
wire net_13534;
wire net_16204;
wire net_15552;
wire net_7162;
wire net_6866;
wire net_3955;
wire net_13770;
wire net_14531;
wire net_16226;
wire net_5950;
wire net_11893;
wire net_8246;
wire net_18852;
wire net_9157;
wire net_18807;
wire net_7252;
wire net_5503;
wire net_2235;
wire net_8303;
wire net_11007;
wire net_11329;
wire net_5846;
wire net_2080;
wire net_3675;
wire net_6714;
wire net_2711;
wire net_18760;
wire net_2097;
wire net_6194;
wire net_11120;
wire net_3619;
wire net_15362;
wire net_1782;
wire net_16828;
wire net_8450;
wire net_11191;
wire net_4863;
wire net_273;
wire net_1278;
wire net_6430;
wire net_4714;
wire net_3182;
wire net_12643;
wire net_2098;
wire net_4232;
wire net_177;
wire net_3355;
wire net_4305;
wire net_18087;
wire net_7806;
wire net_17413;
wire net_8739;
wire net_2803;
wire net_3301;
wire net_6370;
wire net_12133;
wire net_6090;
wire net_17338;
wire net_953;
wire net_17640;
wire net_11600;
wire net_11171;
wire net_1074;
wire net_1058;
wire net_7186;
wire net_12728;
wire net_15911;
wire net_9535;
wire net_11295;
wire net_15954;
wire net_16658;
wire net_6159;
wire x1215;
wire net_9064;
wire net_14004;
wire net_6962;
wire net_2489;
wire net_18063;
wire net_13829;
wire net_3160;
wire net_2125;
wire net_16173;
wire net_7622;
wire net_8179;
wire net_9546;
wire net_13078;
wire net_2623;
wire net_16210;
wire net_261;
wire net_8448;
wire net_17757;
wire net_10654;
wire net_15803;
wire net_2362;
wire net_12837;
wire net_8869;
wire net_18703;
wire net_4456;
wire net_4354;
wire net_5111;
wire net_1955;
wire net_8507;
wire net_8196;
wire net_12886;
wire net_9729;
wire net_18948;
wire net_3012;
wire x13025;
wire net_13134;
wire x27;
wire net_6014;
wire net_5367;
wire net_3754;
wire net_10432;
wire net_17328;
wire net_6075;
wire net_9935;
wire net_18357;
wire net_3989;
wire net_11356;
wire net_13902;
wire net_7304;
wire net_10515;
wire net_5285;
wire net_10875;
wire net_11312;
wire net_1994;
wire net_10499;
wire net_8574;
wire net_4668;
wire net_3897;
wire net_9288;
wire net_17262;
wire net_3960;
wire net_4374;
wire net_15983;
wire net_16732;
wire net_6152;
wire net_3992;
wire net_15959;
wire net_17773;
wire net_2287;
wire net_4211;
wire net_14590;
wire net_18010;
wire net_448;
wire net_8224;
wire net_886;
wire net_3189;
wire net_18466;
wire net_2988;
wire net_18835;
wire net_6811;
wire net_4592;
wire net_16304;
wire net_5279;
wire net_19042;
wire net_3651;
wire net_12182;
wire net_16710;
wire net_9059;
wire net_14345;
wire net_1470;
wire net_11440;
wire net_13358;
wire net_14053;
wire net_4627;
wire net_4423;
wire net_15348;
wire net_14796;
wire net_15373;
wire x13884;
wire net_13674;
wire net_16557;
wire net_4233;
wire net_18090;
wire net_7650;
wire net_4796;
wire x12940;
wire net_15057;
wire net_8289;
wire net_2778;
wire net_13662;
wire net_15148;
wire net_2756;
wire net_12896;
wire net_9605;
wire net_1085;
wire net_592;
wire net_17228;
wire net_9528;
wire net_8983;
wire net_7531;
wire net_2266;
wire net_281;
wire x4607;
wire net_8337;
wire net_12493;
wire net_14699;
wire net_17342;
wire net_5254;
wire net_5193;
wire net_5235;
wire net_16385;
wire net_18143;
wire net_5520;
wire net_15928;
wire net_15344;
wire net_10801;
wire net_10281;
wire net_13532;
wire net_526;
wire net_2718;
wire net_13123;
wire net_2747;
wire net_16331;
wire net_14365;
wire net_18016;
wire net_9232;
wire net_12271;
wire net_16192;
wire net_974;
wire net_12348;
wire net_11777;
wire net_16858;
wire net_923;
wire net_13853;
wire x13069;
wire x3816;
wire net_10947;
wire net_1707;
wire net_4566;
wire net_2190;
wire net_1881;
wire net_7014;
wire net_10487;
wire net_16607;
wire net_10900;
wire net_12925;
wire net_15788;
wire net_3323;
wire net_11697;
wire net_6347;
wire net_7867;
wire net_8961;
wire net_11073;
wire net_12221;
wire net_1492;
wire net_6179;
wire net_14312;
wire net_6363;
wire net_10585;
wire net_9275;
wire net_8267;
wire net_2537;
wire net_11088;
wire net_16966;
wire net_14904;
wire net_18211;
wire net_3767;
wire net_6919;
wire net_6408;
wire net_18773;
wire x13234;
wire net_4105;
wire net_11984;
wire net_11397;
wire net_5594;
wire net_6132;
wire net_9553;
wire net_9193;
wire net_4569;
wire net_5754;
wire net_17379;
wire net_15829;
wire net_17553;
wire net_13000;
wire net_6214;
wire net_9798;
wire net_15944;
wire net_2049;
wire net_2273;
wire net_11558;
wire net_617;
wire net_11026;
wire net_18158;
wire net_6030;
wire net_8656;
wire net_13456;
wire net_4176;
wire net_18486;
wire net_16935;
wire net_18402;
wire net_4032;
wire net_4154;
wire net_17565;
wire net_9294;
wire net_9413;
wire net_9794;
wire net_10420;
wire net_7877;
wire net_9000;
wire net_16505;
wire net_5917;
wire net_5709;
wire net_3870;
wire net_6254;
wire net_18269;
wire net_5456;
wire net_7105;
wire net_15662;
wire net_18383;
wire net_8310;
wire net_5946;
wire net_17296;
wire net_11662;
wire net_16281;
wire net_14481;
wire x13722;
wire net_8742;
wire net_16984;
wire net_6854;
wire net_14132;
wire net_18271;
wire net_12216;
wire net_16560;
wire net_10082;
wire net_13766;
wire net_384;
wire net_4191;
wire net_3503;
wire net_17324;
wire net_17277;
wire net_16051;
wire net_18953;
wire net_5792;
wire net_13366;
wire net_2599;
wire net_15136;
wire x690;
wire net_2665;
wire net_17355;
wire net_3642;
wire net_9200;
wire net_2707;
wire net_7426;
wire net_15834;
wire x4503;
wire net_485;
wire net_11179;
wire net_18106;
wire net_7772;
wire net_15030;
wire net_16394;
wire net_7348;
wire net_11364;
wire net_16669;
wire net_18718;
wire net_11081;
wire net_11589;
wire net_9329;
wire net_13402;
wire net_15822;
wire net_1685;
wire net_4768;
wire x4489;
wire net_17815;
wire net_12019;
wire net_13147;
wire net_14239;
wire net_2644;
wire net_6102;
wire net_12815;
wire net_18862;
wire net_16774;
wire net_13093;
wire net_12686;
wire net_286;
wire net_11668;
wire net_3584;
wire net_7051;
wire net_5588;
wire net_11591;
wire net_4999;
wire net_4340;
wire net_10275;
wire net_4954;
wire net_17971;
wire net_16268;
wire net_5878;
wire net_15588;
wire net_10277;
wire net_3475;
wire net_8423;
wire net_14142;
wire net_5832;
wire net_9070;
wire net_8232;
wire net_1951;
wire net_12608;
wire net_7292;
wire x3561;
wire net_16200;
wire net_12724;
wire net_9759;
wire net_15608;
wire net_8976;
wire net_7661;
wire net_12000;
wire net_15576;
wire net_11869;
wire net_5567;
wire net_2558;
wire net_2040;
wire x4143;
wire net_1508;
wire net_3379;
wire net_931;
wire net_4466;
wire net_18936;
wire net_5983;
wire net_18940;
wire net_2242;
wire net_8505;
wire net_7672;
wire net_6802;
wire net_759;
wire x4840;
wire net_7852;
wire net_11711;
wire net_8832;
wire net_11155;
wire net_8083;
wire net_18376;
wire net_17781;
wire net_6742;
wire net_6428;
wire net_5242;
wire net_17788;
wire net_6924;
wire net_6516;
wire net_12573;
wire net_14585;
wire net_1341;
wire net_17689;
wire net_4541;
wire net_5210;
wire net_3242;
wire net_8138;
wire net_1835;
wire net_18324;
wire net_333;
wire net_15013;
wire net_14491;
wire net_9114;
wire net_9322;
wire net_15203;
wire net_4664;
wire net_15184;
wire net_18333;
wire net_5976;
wire net_13547;
wire net_3923;
wire net_10155;
wire net_8839;
wire net_7210;
wire net_2554;
wire net_16612;
wire net_12196;
wire net_17934;
wire net_4479;
wire net_15708;
wire net_16276;
wire net_7931;
wire net_14453;
wire net_9716;
wire net_14100;
wire net_6354;
wire net_9381;
wire net_13630;
wire net_10928;
wire net_10316;
wire net_7980;
wire net_204;
wire net_14885;
wire net_4596;
wire net_13065;
wire net_12932;
wire x13163;
wire net_14750;
wire net_7626;
wire net_7382;
wire net_16431;
wire net_16402;
wire net_18641;
wire net_14942;
wire net_15461;
wire net_12045;
wire net_15239;
wire net_5416;
wire net_8142;
wire net_17096;
wire net_17161;
wire net_10784;
wire net_1916;
wire net_15941;
wire net_14808;
wire net_11419;
wire net_2468;
wire net_15306;
wire net_7073;
wire net_14416;
wire net_16141;
wire net_10953;
wire net_18412;
wire net_2195;
wire net_11546;
wire net_3421;
wire net_11246;
wire net_1691;
wire net_10089;
wire net_9197;
wire net_18799;
wire net_595;
wire net_12312;
wire net_1320;
wire net_9461;
wire net_9573;
wire net_7434;
wire net_6960;
wire net_8960;
wire net_18050;
wire net_1710;
wire net_10994;
wire net_9017;
wire net_11456;
wire net_14274;
wire net_11922;
wire net_11443;
wire net_15742;
wire net_10524;
wire net_18192;
wire net_18619;
wire net_17625;
wire net_5988;
wire net_6969;
wire net_4336;
wire net_9601;
wire net_13030;
wire net_15699;
wire net_4161;
wire net_3039;
wire net_6207;
wire net_2217;
wire net_938;
wire net_1761;
wire net_12163;
wire net_5682;
wire net_4683;
wire net_183;
wire net_1440;
wire net_7330;
wire net_18424;
wire net_6539;
wire net_1011;
wire net_8792;
wire net_7040;
wire net_1355;
wire net_9902;
wire net_800;
wire net_8420;
wire net_18231;
wire net_9221;
wire net_8847;
wire net_13586;
wire net_18964;
wire net_5992;
wire net_12750;
wire net_11648;
wire net_4046;
wire net_9405;
wire net_16733;
wire net_2580;
wire net_13834;
wire net_9696;
wire net_13997;
wire x13514;
wire net_15994;
wire net_1643;
wire net_1385;
wire net_9961;
wire net_13302;
wire net_1534;
wire net_1919;
wire net_15029;
wire net_9836;
wire net_19007;
wire net_12843;
wire net_8992;
wire net_14162;
wire net_4876;
wire net_18566;
wire net_16234;
wire net_659;
wire net_9087;
wire net_14860;
wire net_8993;
wire net_14652;
wire net_899;
wire net_1010;
wire net_10224;
wire net_18873;
wire net_3654;
wire net_13883;
wire net_10139;
wire net_15542;
wire net_15082;
wire net_18579;
wire net_2908;
wire net_14830;
wire net_4981;
wire x43;
wire net_14566;
wire net_15020;
wire net_16083;
wire net_13594;
wire net_13780;
wire net_14576;
wire net_13813;
wire net_4449;
wire net_16720;
wire net_7339;
wire net_6458;
wire net_11929;
wire net_2675;
wire net_2794;
wire net_13528;
wire net_13567;
wire net_6986;
wire net_16633;
wire net_1752;
wire net_2527;
wire net_11906;
wire net_2091;
wire net_14478;
wire net_17594;
wire net_2406;
wire net_6289;
wire net_8722;
wire net_17157;
wire net_18397;
wire net_807;
wire net_3405;
wire net_3270;
wire net_12422;
wire net_15456;
wire net_12665;
wire net_6880;
wire net_10238;
wire net_2474;
wire net_13931;
wire net_2530;
wire net_11578;
wire net_15824;
wire net_9472;
wire net_6192;
wire net_217;
wire net_7679;
wire net_18070;
wire net_14935;
wire net_5336;
wire net_12086;
wire net_915;
wire net_8844;
wire net_5634;
wire net_2226;
wire net_3849;
wire net_17016;
wire net_8099;
wire net_8909;
wire net_18637;
wire net_8028;
wire net_17306;
wire net_14700;
wire net_15479;
wire net_8369;
wire net_2863;
wire net_3507;
wire net_1165;
wire net_5167;
wire net_677;
wire net_1472;
wire net_18727;
wire net_2939;
wire net_1113;
wire net_13294;
wire net_9945;
wire net_17894;
wire net_11208;
wire net_11619;
wire net_15316;
wire net_18442;
wire net_7464;
wire net_8362;
wire net_11040;
wire net_5120;
wire net_15197;
wire net_14969;
wire net_5948;
wire net_5676;
wire net_15484;
wire net_8357;
wire net_2658;
wire net_2174;
wire net_14875;
wire net_784;
wire net_16460;
wire net_8481;
wire net_8751;
wire net_6021;
wire net_18173;
wire net_2326;
wire x1804;
wire net_11566;
wire net_3540;
wire net_8094;
wire net_11234;
wire net_5375;
wire net_9489;
wire net_18431;
wire net_12078;
wire net_19036;
wire net_17125;
wire net_1318;
wire net_3238;
wire net_10677;
wire net_15227;
wire net_15486;
wire net_16480;
wire net_7155;
wire net_4349;
wire net_3575;
wire net_11195;
wire net_8023;
wire net_18240;
wire net_6440;
wire net_15039;
wire net_4984;
wire net_306;
wire net_18127;
wire net_4516;
wire net_5371;
wire net_9026;
wire net_5061;
wire net_6471;
wire net_2610;
wire net_4432;
wire net_4584;
wire net_1329;
wire net_14391;
wire net_362;
wire net_3127;
wire net_9959;
wire net_1052;
wire net_3831;
wire net_11180;
wire net_13974;
wire net_18163;
wire net_9477;
wire net_17966;
wire net_17004;
wire net_15083;
wire net_4859;
wire net_6413;
wire net_226;
wire net_18856;
wire net_18367;
wire net_7015;
wire net_9160;
wire net_16169;
wire net_2887;
wire net_4207;
wire net_15515;
wire net_7741;
wire net_1983;
wire net_8735;
wire net_10129;
wire net_10248;
wire net_3030;
wire net_10251;
wire net_3842;
wire net_15433;
wire net_4266;
wire net_1553;
wire net_13421;
wire net_2491;
wire net_8819;
wire net_10563;
wire net_3208;
wire net_2704;
wire net_10933;
wire net_15591;
wire net_5819;
wire net_14663;
wire net_3910;
wire net_1851;
wire net_13684;
wire net_3445;
wire net_10976;
wire net_18470;
wire net_8709;
wire net_2941;
wire net_477;
wire net_3348;
wire x13134;
wire net_17368;
wire net_2943;
wire net_9377;
wire net_3861;
wire net_10892;
wire net_6758;
wire net_6905;
wire net_2315;
wire net_8325;
wire net_2231;
wire net_15501;
wire net_17582;
wire net_14646;
wire net_3812;
wire net_1200;
wire net_9595;
wire net_17136;
wire net_9509;
wire net_18429;
wire net_12329;
wire net_7558;
wire net_11135;
wire net_11487;
wire net_13980;
wire net_16675;
wire net_3437;
wire net_18391;
wire net_19024;
wire net_472;
wire net_1510;
wire net_14286;
wire net_14022;
wire net_3077;
wire net_18401;
wire net_8639;
wire net_4829;
wire net_13608;
wire net_9430;
wire net_4171;
wire net_1528;
wire net_12676;
wire net_13579;
wire net_15628;
wire net_1749;
wire net_3367;
wire net_4915;
wire x2451;
wire net_4784;
wire net_8386;
wire net_12355;
wire net_601;
wire net_1362;
wire net_4385;
wire net_2346;
wire net_829;
wire net_9315;
wire net_13025;
wire net_12396;
wire net_2294;
wire net_11856;
wire net_13867;
wire net_4978;
wire net_14174;
wire net_2393;
wire net_18646;
wire net_3917;
wire net_15171;
wire net_8539;
wire net_8812;
wire net_3376;
wire net_13671;
wire net_7979;
wire net_16351;
wire net_13845;
wire net_14926;
wire net_15090;
wire net_17983;
wire net_17174;
wire net_7218;
wire net_5319;
wire net_11045;
wire net_6357;
wire net_3750;
wire net_12637;
wire net_5314;
wire net_5749;
wire net_2696;
wire net_9687;
wire net_10464;
wire net_12736;
wire net_6026;
wire net_14168;
wire net_8457;
wire net_10457;
wire net_1449;
wire net_16222;
wire net_6984;
wire net_5618;
wire x13464;
wire net_15740;
wire net_5310;
wire net_9725;
wire net_8620;
wire net_13114;
wire net_1220;
wire net_12989;
wire net_14729;
wire net_17420;
wire net_12343;
wire net_4693;
wire net_4017;
wire net_11394;
wire net_10194;
wire net_6346;
wire net_12716;
wire net_11781;
wire net_4945;
wire net_18046;
wire net_15097;
wire net_14208;
wire net_2334;
wire net_17213;
wire net_1367;
wire net_7943;
wire net_16644;
wire net_17531;
wire net_7960;
wire net_18817;
wire net_4079;
wire x13185;
wire net_12104;
wire net_1371;
wire net_12542;
wire net_13511;
wire net_16769;
wire net_5002;
wire net_8054;
wire net_18441;
wire net_6609;
wire net_7837;
wire net_16420;
wire net_16261;
wire net_6517;
wire net_4704;
wire net_15526;
wire net_5782;
wire net_9843;
wire net_7864;
wire net_11885;
wire net_10359;
wire net_11826;
wire net_1461;
wire net_18008;
wire net_17859;
wire net_12799;
wire net_7512;
wire net_16762;
wire net_3177;
wire net_15769;
wire net_8270;
wire net_11325;
wire net_10011;
wire net_12556;
wire net_14526;
wire net_7222;
wire net_9459;
wire net_15921;
wire net_8891;
wire x3803;
wire x3762;
wire net_10360;
wire net_10475;
wire net_437;
wire net_10568;
wire net_3573;
wire net_13208;
wire net_16926;
wire net_9861;
wire net_10390;
wire net_11477;
wire net_7371;
wire net_9071;
wire net_10855;
wire net_12498;
wire net_7140;
wire net_17113;
wire net_624;
wire net_2148;
wire net_15669;
wire net_11616;
wire net_14427;
wire net_16295;
wire net_8517;
wire net_14063;
wire net_6005;
wire net_688;
wire net_8732;
wire x1340;
wire net_5808;
wire net_8170;
wire net_3027;
wire net_12777;
wire net_16927;
wire net_17912;
wire net_5343;
wire net_14464;
wire net_6625;
wire net_15659;
wire net_15999;
wire net_9940;
wire net_15813;
wire net_5497;
wire net_4096;
wire net_7924;
wire net_16587;
wire net_5214;
wire net_4822;
wire net_3986;
wire x771;
wire net_11754;
wire net_7482;
wire net_1243;
wire net_6839;
wire net_1660;
wire net_12035;
wire net_1484;
wire net_5864;
wire net_3667;
wire net_6566;
wire net_9949;
wire net_6041;
wire net_1635;
wire net_6779;
wire net_5027;
wire net_4840;
wire net_12697;
wire net_7133;
wire net_7523;
wire net_8828;
wire net_7174;
wire net_6871;
wire net_10306;
wire net_7020;
wire net_3002;
wire net_16241;
wire net_854;
wire net_17850;
wire net_2619;
wire net_8713;
wire net_5559;
wire net_18351;
wire net_2221;
wire net_15585;
wire net_11424;
wire net_6959;
wire net_5264;
wire net_10369;
wire net_6447;
wire net_7789;
wire net_18606;
wire net_16873;
wire net_18625;
wire x154;
wire net_9181;
wire net_5746;
wire net_16366;
wire net_4643;
wire net_332;
wire net_1745;
wire net_13601;
wire net_1679;
wire net_7364;
wire net_4883;
wire net_9058;
wire net_13739;
wire net_656;
wire net_5723;
wire net_4800;
wire net_8489;
wire net_18371;
wire net_17180;
wire net_8935;
wire net_4284;
wire net_7027;
wire net_16316;
wire net_3113;
wire net_17033;
wire net_10924;
wire net_14157;
wire net_8826;
wire net_6816;
wire net_8614;
wire net_15974;
wire net_3969;
wire net_7232;
wire net_13266;
wire net_14768;
wire net_6602;
wire net_9873;
wire net_11164;
wire net_12615;
wire net_7688;
wire net_17732;
wire net_15198;
wire net_6162;
wire net_17765;
wire net_1698;
wire net_5897;
wire net_18756;
wire net_1017;
wire net_12391;
wire net_14309;
wire net_14379;
wire net_18722;
wire net_13334;
wire net_14293;
wire net_412;
wire net_4798;
wire net_8887;
wire net_16090;
wire net_9869;
wire net_1873;
wire net_3801;
wire net_453;
wire net_7547;
wire net_10209;
wire net_17139;
wire net_5835;
wire net_18450;
wire net_2263;
wire net_10439;
wire net_6181;
wire net_3624;
wire net_7967;
wire net_9391;
wire x963;
wire net_951;
wire net_2086;
wire net_11596;
wire net_17382;
wire net_4930;
wire net_18665;
wire net_17252;
wire net_16715;
wire net_12278;
wire net_12869;
wire net_7272;
wire net_7096;
wire net_8977;
wire net_12654;
wire net_18517;
wire net_10222;
wire net_14389;
wire net_10648;
wire net_12350;
wire net_12121;
wire net_2966;
wire net_15146;
wire net_1253;
wire net_13186;
wire net_2500;
wire net_9808;
wire net_10508;
wire net_17716;
wire net_13971;
wire net_3900;
wire net_13315;
wire x13414;
wire net_15889;
wire net_3153;
wire net_16456;
wire net_6721;
wire net_5471;
wire net_5155;
wire x13145;
wire net_3598;
wire net_16418;
wire net_3938;
wire net_8676;
wire net_7534;
wire x12915;
wire net_11289;
wire net_15757;
wire net_9592;
wire net_18669;
wire net_1502;
wire net_11282;
wire net_6596;
wire net_11065;
wire net_10329;
wire net_11306;
wire net_640;
wire net_10117;
wire net_12138;
wire net_7508;
wire net_775;
wire net_752;
wire net_10903;
wire net_18114;
wire net_498;
wire net_535;
wire net_3716;
wire net_17387;
wire net_2721;
wire net_8900;
wire net_2637;
wire net_15380;
wire net_6768;
wire net_4902;
wire net_5419;
wire net_299;
wire net_12228;
wire net_18266;
wire net_12894;
wire net_7413;
wire net_12387;
wire net_2024;
wire net_11755;
wire net_3254;
wire net_11549;
wire net_9569;
wire net_9779;
wire net_9040;
wire net_3725;
wire net_17809;
wire net_15569;
wire net_9111;
wire net_6088;
wire net_5857;
wire net_5041;
wire net_15161;
wire net_407;
wire net_4405;
wire net_16903;
wire net_11793;
wire net_18884;
wire net_8723;
wire net_9801;
wire net_2312;
wire net_16547;
wire net_8586;
wire net_2073;
wire net_8189;
wire net_9146;
wire net_4057;
wire net_5105;
wire net_14244;
wire net_6081;
wire net_14975;
wire net_14863;
wire net_16374;
wire net_5507;
wire net_12173;
wire net_12526;
wire net_7565;
wire net_15339;
wire net_1981;
wire net_4302;
wire net_6245;
wire net_1218;
wire net_10606;
wire net_15042;
wire net_16128;
wire net_3286;
wire net_11430;
wire net_15604;
wire net_1398;
wire x1152;
wire net_12432;
wire net_13219;
wire net_10503;
wire net_4399;
wire net_8197;
wire net_6117;
wire net_1144;
wire net_8297;
wire net_16373;
wire net_17571;
wire net_10646;
wire net_2260;
wire net_2865;
wire net_3606;
wire net_9770;
wire net_17116;
wire net_702;
wire net_4328;
wire net_1477;
wire net_3195;
wire net_3210;
wire net_16013;
wire net_3318;
wire net_13221;
wire net_7800;
wire net_8188;
wire net_17674;
wire net_8122;
wire net_7571;
wire net_11682;
wire net_12948;
wire net_12904;
wire net_15214;
wire net_1193;
wire net_12979;
wire net_9412;
wire net_1425;
wire net_17331;
wire net_17068;
wire net_8436;
wire net_10790;
wire net_1813;
wire net_10622;
wire net_18406;
wire net_10673;
wire net_7945;
wire net_17363;
wire net_12411;
wire net_983;
wire net_18992;
wire net_16651;
wire net_355;
wire net_7258;
wire net_13702;
wire net_9513;
wire net_8102;
wire net_12427;
wire net_15534;
wire net_7311;
wire net_723;
wire net_11341;
wire net_7614;
wire net_2483;
wire net_18068;
wire net_16080;
wire net_12026;
wire net_14608;
wire net_10202;
wire net_10501;
wire net_15096;
wire net_10547;
wire net_19013;
wire net_16388;
wire net_3948;
wire net_6142;
wire net_13475;
wire net_13455;
wire net_12414;
wire net_12872;
wire net_9493;
wire net_8254;
wire net_11945;
wire net_3819;
wire net_15640;
wire net_254;
wire net_1501;
wire net_3003;
wire net_12103;
wire net_574;
wire net_11375;

// Start cells
SDFF_X2 inst_1783 ( .D(net_7291), .SI(net_6908), .Q(net_6908), .SE(net_6284), .CK(net_15340) );
CLKBUF_X2 inst_17321 ( .A(net_17168), .Z(net_17169) );
CLKBUF_X2 inst_18950 ( .A(net_18797), .Z(net_18798) );
CLKBUF_X2 inst_17160 ( .A(net_17007), .Z(net_17008) );
SDFFR_X1 inst_2685 ( .SI(net_7547), .SE(net_5043), .CK(net_9684), .RN(x6501), .Q(x3968), .D(x3968) );
INV_X4 inst_5359 ( .A(net_1465), .ZN(net_1145) );
CLKBUF_X2 inst_16895 ( .A(net_16742), .Z(net_16743) );
CLKBUF_X2 inst_13828 ( .A(net_13675), .Z(net_13676) );
INV_X2 inst_6439 ( .A(net_1273), .ZN(net_640) );
INV_X4 inst_5306 ( .ZN(net_1704), .A(net_1478) );
SDFFR_X2 inst_2205 ( .Q(net_7448), .D(net_7448), .SE(net_2863), .CK(net_12825), .SI(x13594), .RN(x6501) );
CLKBUF_X2 inst_17222 ( .A(net_16127), .Z(net_17070) );
OR2_X4 inst_2858 ( .A1(net_6808), .A2(net_6805), .ZN(net_613) );
AOI21_X2 inst_8981 ( .ZN(net_1934), .A(net_1933), .B1(net_1756), .B2(net_1755) );
INV_X4 inst_5488 ( .ZN(net_1267), .A(net_726) );
CLKBUF_X2 inst_19173 ( .A(net_15886), .Z(net_19021) );
CLKBUF_X2 inst_13926 ( .A(net_13773), .Z(net_13774) );
CLKBUF_X2 inst_15089 ( .A(net_14182), .Z(net_14937) );
XNOR2_X2 inst_214 ( .ZN(net_1447), .B(net_1446), .A(net_1269) );
CLKBUF_X2 inst_13990 ( .A(net_13837), .Z(net_13838) );
CLKBUF_X2 inst_18233 ( .A(net_18080), .Z(net_18081) );
CLKBUF_X2 inst_15915 ( .A(net_11494), .Z(net_15763) );
AND2_X4 inst_9115 ( .ZN(net_1740), .A2(net_1260), .A1(net_1259) );
SDFF_X2 inst_548 ( .Q(net_8693), .D(net_8693), .SI(net_3975), .SE(net_3935), .CK(net_10272) );
CLKBUF_X2 inst_16093 ( .A(net_15940), .Z(net_15941) );
NAND2_X2 inst_4372 ( .A1(net_7114), .A2(net_5164), .ZN(net_5085) );
CLKBUF_X2 inst_18084 ( .A(net_17931), .Z(net_17932) );
DFFR_X2 inst_7191 ( .QN(net_8955), .D(net_2422), .CK(net_15064), .RN(x6501) );
CLKBUF_X2 inst_12796 ( .A(net_12643), .Z(net_12644) );
CLKBUF_X2 inst_14747 ( .A(net_14594), .Z(net_14595) );
AOI22_X2 inst_8488 ( .B1(net_6545), .A1(net_6512), .A2(net_6137), .B2(net_6104), .ZN(net_3452) );
CLKBUF_X2 inst_14178 ( .A(net_14025), .Z(net_14026) );
CLKBUF_X2 inst_17516 ( .A(net_17363), .Z(net_17364) );
CLKBUF_X2 inst_14148 ( .A(net_13995), .Z(net_13996) );
CLKBUF_X2 inst_13127 ( .A(net_10097), .Z(net_12975) );
INV_X2 inst_6406 ( .ZN(net_1073), .A(net_1072) );
CLKBUF_X2 inst_18400 ( .A(net_18247), .Z(net_18248) );
CLKBUF_X2 inst_12400 ( .A(net_12247), .Z(net_12248) );
SDFF_X2 inst_1228 ( .Q(net_7954), .D(net_7954), .SE(net_2755), .SI(net_2574), .CK(net_16086) );
AOI21_X2 inst_8913 ( .ZN(net_5805), .A(net_5745), .B2(net_5607), .B1(net_5256) );
CLKBUF_X2 inst_13185 ( .A(net_11608), .Z(net_13033) );
NAND2_X2 inst_4221 ( .A1(net_6894), .A2(net_5247), .ZN(net_5239) );
SDFF_X2 inst_521 ( .Q(net_8876), .D(net_8876), .SI(net_3955), .SE(net_3936), .CK(net_11017) );
INV_X2 inst_6534 ( .A(net_6467), .ZN(net_520) );
INV_X4 inst_5947 ( .A(net_8971), .ZN(net_524) );
NAND2_X2 inst_4473 ( .A2(net_5657), .ZN(net_4644), .A1(net_2697) );
SDFF_X2 inst_1685 ( .SI(net_7721), .Q(net_7721), .D(net_2719), .SE(net_2559), .CK(net_18767) );
SDFFR_X2 inst_2511 ( .Q(net_8997), .D(net_8997), .SI(net_2632), .SE(net_2562), .CK(net_14524), .RN(x6501) );
CLKBUF_X2 inst_12320 ( .A(net_10751), .Z(net_12168) );
AND4_X2 inst_9038 ( .A4(net_1819), .ZN(net_1649), .A2(net_1648), .A1(net_1501), .A3(net_587) );
DFFS_X2 inst_6910 ( .QN(net_7209), .D(net_2255), .CK(net_15174), .SN(x6501) );
NOR2_X2 inst_3578 ( .A2(net_9057), .A1(net_9054), .ZN(net_1458) );
CLKBUF_X2 inst_9257 ( .A(net_9104), .Z(net_9105) );
CLKBUF_X2 inst_15477 ( .A(net_15324), .Z(net_15325) );
CLKBUF_X2 inst_14731 ( .A(net_14578), .Z(net_14579) );
CLKBUF_X2 inst_9938 ( .A(net_9785), .Z(net_9786) );
CLKBUF_X2 inst_12238 ( .A(net_12085), .Z(net_12086) );
INV_X4 inst_5940 ( .A(net_7244), .ZN(net_1942) );
CLKBUF_X2 inst_17892 ( .A(net_15610), .Z(net_17740) );
CLKBUF_X2 inst_18107 ( .A(net_11159), .Z(net_17955) );
CLKBUF_X2 inst_14010 ( .A(net_13857), .Z(net_13858) );
CLKBUF_X2 inst_13236 ( .A(net_9598), .Z(net_13084) );
CLKBUF_X2 inst_10825 ( .A(net_10672), .Z(net_10673) );
NOR2_X2 inst_3392 ( .ZN(net_4640), .A2(net_4473), .A1(net_4412) );
CLKBUF_X2 inst_18376 ( .A(net_18223), .Z(net_18224) );
INV_X2 inst_6232 ( .ZN(net_5478), .A(net_5298) );
SDFFR_X2 inst_2342 ( .SE(net_2260), .Q(net_364), .D(net_364), .CK(net_11458), .RN(x6501), .SI(x1829) );
CLKBUF_X2 inst_15849 ( .A(net_15696), .Z(net_15697) );
AND2_X4 inst_9143 ( .A2(net_8948), .A1(net_6113), .ZN(net_1324) );
SDFF_X2 inst_1617 ( .Q(net_8159), .D(net_8159), .SI(net_2720), .SE(net_2538), .CK(net_18373) );
CLKBUF_X2 inst_12553 ( .A(net_10760), .Z(net_12401) );
XNOR2_X2 inst_151 ( .ZN(net_2040), .B(net_2039), .A(net_1933) );
SDFFR_X2 inst_2256 ( .D(net_7387), .SE(net_2797), .SI(net_196), .Q(net_196), .CK(net_14766), .RN(x6501) );
CLKBUF_X2 inst_18916 ( .A(net_18763), .Z(net_18764) );
DFFR_X1 inst_7519 ( .Q(net_340), .D(net_298), .CK(net_16164), .RN(x6501) );
NAND2_X2 inst_4880 ( .A1(net_8280), .ZN(net_782), .A2(net_488) );
CLKBUF_X2 inst_11637 ( .A(net_11484), .Z(net_11485) );
CLKBUF_X2 inst_10370 ( .A(net_10217), .Z(net_10218) );
NAND3_X4 inst_3867 ( .A3(net_6261), .A1(net_6191), .ZN(net_4817), .A2(net_4816) );
SDFFS_X2 inst_2072 ( .SI(net_7388), .SE(net_2795), .Q(net_177), .D(net_177), .CK(net_17435), .SN(x6501) );
SDFF_X2 inst_1603 ( .Q(net_8139), .D(net_8139), .SI(net_2639), .SE(net_2541), .CK(net_16484) );
CLKBUF_X2 inst_9634 ( .A(net_9084), .Z(net_9482) );
SDFF_X2 inst_340 ( .SI(net_8610), .Q(net_8610), .SE(net_3984), .D(net_3967), .CK(net_13073) );
CLKBUF_X2 inst_18322 ( .A(net_18169), .Z(net_18170) );
CLKBUF_X2 inst_14978 ( .A(net_14825), .Z(net_14826) );
AOI22_X2 inst_8109 ( .B1(net_7941), .A1(net_7839), .B2(net_6103), .A2(net_4398), .ZN(net_4038) );
CLKBUF_X2 inst_11075 ( .A(net_10922), .Z(net_10923) );
NAND2_X2 inst_4280 ( .A1(net_7005), .A2(net_5249), .ZN(net_5180) );
AOI22_X2 inst_8171 ( .B1(net_8566), .A1(net_8455), .A2(net_6263), .B2(net_6262), .ZN(net_3859) );
DFFR_X1 inst_7493 ( .D(net_3213), .CK(net_14515), .RN(x6501), .Q(x933) );
INV_X4 inst_5411 ( .ZN(net_2408), .A(net_872) );
CLKBUF_X2 inst_18543 ( .A(net_18390), .Z(net_18391) );
CLKBUF_X2 inst_14279 ( .A(net_14126), .Z(net_14127) );
NAND2_X2 inst_4244 ( .A1(net_7025), .A2(net_5249), .ZN(net_5216) );
SDFF_X2 inst_1490 ( .SI(net_7263), .Q(net_7040), .D(net_7040), .SE(net_6280), .CK(net_17072) );
CLKBUF_X2 inst_15421 ( .A(net_9059), .Z(net_15269) );
NAND2_X2 inst_4559 ( .ZN(net_3888), .A2(net_3887), .A1(net_3251) );
NAND4_X2 inst_3709 ( .ZN(net_4428), .A4(net_4334), .A1(net_3707), .A2(net_3706), .A3(net_3705) );
CLKBUF_X2 inst_10934 ( .A(net_10781), .Z(net_10782) );
INV_X2 inst_6319 ( .ZN(net_3344), .A(net_3289) );
SDFF_X2 inst_827 ( .SI(net_8487), .Q(net_8487), .D(net_3965), .SE(net_3884), .CK(net_13030) );
CLKBUF_X2 inst_18560 ( .A(net_18407), .Z(net_18408) );
CLKBUF_X2 inst_15309 ( .A(net_11274), .Z(net_15157) );
CLKBUF_X2 inst_11477 ( .A(net_11324), .Z(net_11325) );
CLKBUF_X2 inst_17498 ( .A(net_17345), .Z(net_17346) );
CLKBUF_X2 inst_9573 ( .A(net_9420), .Z(net_9421) );
CLKBUF_X2 inst_15231 ( .A(net_15078), .Z(net_15079) );
CLKBUF_X2 inst_10730 ( .A(net_9770), .Z(net_10578) );
CLKBUF_X2 inst_10574 ( .A(net_10421), .Z(net_10422) );
DFFR_X2 inst_7140 ( .QN(net_7211), .D(net_2942), .CK(net_15208), .RN(x6501) );
OAI21_X2 inst_3040 ( .B2(net_8235), .B1(net_4928), .ZN(net_4830), .A(net_3273) );
CLKBUF_X2 inst_12937 ( .A(net_12784), .Z(net_12785) );
NAND3_X4 inst_3870 ( .A1(net_6275), .A2(net_6261), .ZN(net_4813), .A3(net_4708) );
CLKBUF_X2 inst_16707 ( .A(net_12525), .Z(net_16555) );
INV_X4 inst_5675 ( .A(net_7606), .ZN(net_2139) );
CLKBUF_X2 inst_17052 ( .A(net_16866), .Z(net_16900) );
NAND2_X2 inst_4640 ( .ZN(net_2797), .A2(net_2418), .A1(net_2116) );
XOR2_X2 inst_18 ( .Z(net_1420), .B(net_1419), .A(net_603) );
INV_X4 inst_6047 ( .A(net_7398), .ZN(net_499) );
NAND2_X2 inst_4128 ( .ZN(net_5396), .A1(net_5128), .A2(net_5127) );
AND3_X4 inst_9040 ( .ZN(net_4362), .A1(net_2644), .A2(net_1803), .A3(net_1624) );
CLKBUF_X2 inst_10154 ( .A(net_9609), .Z(net_10002) );
NAND2_X2 inst_4861 ( .ZN(net_1511), .A2(net_850), .A1(net_180) );
INV_X4 inst_5183 ( .ZN(net_2826), .A(net_2759) );
NAND3_X2 inst_3936 ( .ZN(net_4941), .A3(net_4707), .A1(net_4703), .A2(net_4646) );
CLKBUF_X2 inst_13738 ( .A(net_13585), .Z(net_13586) );
CLKBUF_X2 inst_17866 ( .A(net_15063), .Z(net_17714) );
INV_X4 inst_6069 ( .A(net_6286), .ZN(net_2668) );
CLKBUF_X2 inst_17612 ( .A(net_17459), .Z(net_17460) );
HA_X1 inst_6675 ( .S(net_3166), .CO(net_3165), .B(net_2980), .A(x2400) );
INV_X4 inst_6020 ( .A(net_7647), .ZN(net_667) );
CLKBUF_X2 inst_12739 ( .A(net_12586), .Z(net_12587) );
CLKBUF_X2 inst_14663 ( .A(net_14510), .Z(net_14511) );
CLKBUF_X2 inst_9217 ( .A(net_9060), .Z(net_9065) );
INV_X2 inst_6475 ( .ZN(net_850), .A(net_224) );
DFFR_X2 inst_7364 ( .Q(net_7325), .CK(net_11755), .D(x13047), .RN(x6501) );
INV_X4 inst_5816 ( .A(net_6486), .ZN(net_2876) );
CLKBUF_X2 inst_18259 ( .A(net_16870), .Z(net_18107) );
SDFFR_X1 inst_2695 ( .SI(net_7557), .SE(net_5043), .CK(net_12727), .RN(x6501), .Q(x3816), .D(x3816) );
CLKBUF_X2 inst_13801 ( .A(net_13648), .Z(net_13649) );
CLKBUF_X2 inst_18158 ( .A(net_10437), .Z(net_18006) );
CLKBUF_X2 inst_14833 ( .A(net_14680), .Z(net_14681) );
CLKBUF_X2 inst_12515 ( .A(net_9465), .Z(net_12363) );
CLKBUF_X2 inst_13635 ( .A(net_13482), .Z(net_13483) );
CLKBUF_X2 inst_14980 ( .A(net_14827), .Z(net_14828) );
CLKBUF_X2 inst_10692 ( .A(net_10539), .Z(net_10540) );
CLKBUF_X2 inst_14150 ( .A(net_13997), .Z(net_13998) );
CLKBUF_X2 inst_13228 ( .A(net_13075), .Z(net_13076) );
NOR2_X2 inst_3521 ( .A2(net_3023), .ZN(net_1731), .A1(net_1188) );
AOI21_X2 inst_8969 ( .B2(net_2963), .ZN(net_2914), .B1(net_2913), .A(net_2783) );
NOR2_X2 inst_3440 ( .A2(net_3093), .ZN(net_3055), .A1(net_2815) );
INV_X4 inst_5802 ( .A(net_7224), .ZN(net_2931) );
NAND3_X2 inst_4001 ( .A1(net_7214), .A3(net_7212), .ZN(net_3162), .A2(net_602) );
CLKBUF_X2 inst_12249 ( .A(net_12096), .Z(net_12097) );
AOI22_X2 inst_7897 ( .B1(net_8980), .A2(net_5538), .B2(net_5456), .ZN(net_4532), .A1(net_409) );
AND2_X2 inst_9188 ( .ZN(net_1948), .A1(net_1762), .A2(net_1761) );
INV_X2 inst_6184 ( .ZN(net_5837), .A(net_5781) );
CLKBUF_X2 inst_10958 ( .A(net_10524), .Z(net_10806) );
CLKBUF_X2 inst_18869 ( .A(net_17395), .Z(net_18717) );
CLKBUF_X2 inst_14388 ( .A(net_14235), .Z(net_14236) );
CLKBUF_X2 inst_14922 ( .A(net_14769), .Z(net_14770) );
CLKBUF_X2 inst_10106 ( .A(net_9953), .Z(net_9954) );
SDFF_X2 inst_1027 ( .SI(net_7310), .Q(net_6750), .D(net_6750), .SE(net_3124), .CK(net_11900) );
AOI22_X2 inst_8432 ( .B1(net_6532), .A1(net_6499), .A2(net_6137), .B2(net_6104), .ZN(net_3509) );
SDFF_X2 inst_1143 ( .SI(net_7322), .Q(net_6597), .D(net_6597), .SE(net_3069), .CK(net_11367) );
CLKBUF_X2 inst_11336 ( .A(net_11091), .Z(net_11184) );
CLKBUF_X2 inst_12024 ( .A(net_11126), .Z(net_11872) );
CLKBUF_X2 inst_10457 ( .A(net_10304), .Z(net_10305) );
CLKBUF_X2 inst_12679 ( .A(net_10804), .Z(net_12527) );
CLKBUF_X2 inst_11824 ( .A(net_10877), .Z(net_11672) );
AOI22_X2 inst_8503 ( .B1(net_6615), .A1(net_6582), .A2(net_6257), .B2(net_6110), .ZN(net_3437) );
CLKBUF_X2 inst_18874 ( .A(net_18721), .Z(net_18722) );
NAND2_X2 inst_4147 ( .ZN(net_5371), .A2(net_5212), .A1(net_5108) );
SDFF_X2 inst_1538 ( .Q(net_7991), .D(net_7991), .SI(net_2576), .SE(net_2542), .CK(net_16051) );
CLKBUF_X2 inst_15273 ( .A(net_15120), .Z(net_15121) );
CLKBUF_X2 inst_10349 ( .A(net_10196), .Z(net_10197) );
CLKBUF_X2 inst_12525 ( .A(net_11734), .Z(net_12373) );
INV_X2 inst_6465 ( .A(net_6353), .ZN(net_2145) );
INV_X2 inst_6312 ( .ZN(net_3892), .A(net_3589) );
SDFFR_X2 inst_2179 ( .QN(net_7564), .D(net_3977), .SE(net_3144), .SI(net_3108), .CK(net_10787), .RN(x6501) );
SDFFR_X2 inst_2578 ( .D(net_7394), .QN(net_7254), .SI(net_1958), .SE(net_1379), .CK(net_15352), .RN(x6501) );
DFFR_X1 inst_7514 ( .D(net_7629), .QN(net_7620), .CK(net_15717), .RN(x6501) );
SDFF_X2 inst_1996 ( .SI(net_7921), .Q(net_7921), .D(net_2720), .SE(net_2461), .CK(net_18024) );
CLKBUF_X2 inst_12838 ( .A(net_12685), .Z(net_12686) );
NOR2_X4 inst_3340 ( .A1(net_6141), .A2(net_6140), .ZN(net_1097) );
NAND2_X2 inst_4683 ( .ZN(net_2234), .A1(net_600), .A2(net_265) );
CLKBUF_X2 inst_17414 ( .A(net_17261), .Z(net_17262) );
SDFF_X2 inst_1380 ( .Q(net_8153), .D(net_8153), .SI(net_2658), .SE(net_2538), .CK(net_15290) );
CLKBUF_X2 inst_15890 ( .A(net_15737), .Z(net_15738) );
NAND3_X2 inst_3891 ( .ZN(net_5647), .A1(net_5576), .A3(net_5510), .A2(net_5430) );
CLKBUF_X2 inst_11298 ( .A(net_10122), .Z(net_11146) );
CLKBUF_X2 inst_12484 ( .A(net_12331), .Z(net_12332) );
AOI22_X2 inst_8318 ( .B1(net_8854), .A1(net_8299), .B2(net_6252), .A2(net_4345), .ZN(net_3727) );
CLKBUF_X2 inst_17924 ( .A(net_17771), .Z(net_17772) );
NAND2_X2 inst_4834 ( .A1(net_8903), .ZN(net_1371), .A2(net_1028) );
NOR2_X2 inst_3472 ( .ZN(net_2437), .A2(net_2281), .A1(net_1719) );
AOI221_X4 inst_8736 ( .B1(net_8819), .C1(net_8338), .C2(net_6265), .B2(net_6253), .ZN(net_4330), .A(net_4236) );
CLKBUF_X2 inst_9933 ( .A(net_9780), .Z(net_9781) );
SDFFR_X2 inst_2322 ( .SE(net_2260), .Q(net_352), .D(net_352), .CK(net_11470), .RN(x6501), .SI(x2195) );
SDFF_X2 inst_513 ( .Q(net_8866), .D(net_8866), .SI(net_3959), .SE(net_3936), .CK(net_13203) );
CLKBUF_X2 inst_17725 ( .A(net_17572), .Z(net_17573) );
CLKBUF_X2 inst_14340 ( .A(net_14187), .Z(net_14188) );
SDFF_X2 inst_1630 ( .Q(net_8175), .D(net_8175), .SI(net_2660), .SE(net_2538), .CK(net_17067) );
SDFF_X2 inst_1586 ( .Q(net_8042), .D(net_8042), .SI(net_2656), .SE(net_2545), .CK(net_16717) );
CLKBUF_X2 inst_16624 ( .A(net_16471), .Z(net_16472) );
CLKBUF_X2 inst_9318 ( .A(net_9061), .Z(net_9166) );
CLKBUF_X2 inst_18584 ( .A(net_18431), .Z(net_18432) );
CLKBUF_X2 inst_13954 ( .A(net_13801), .Z(net_13802) );
INV_X4 inst_6083 ( .A(net_6307), .ZN(net_2684) );
NAND2_X2 inst_4256 ( .A1(net_7030), .A2(net_5249), .ZN(net_5204) );
CLKBUF_X2 inst_18416 ( .A(net_9329), .Z(net_18264) );
CLKBUF_X2 inst_10773 ( .A(net_10620), .Z(net_10621) );
CLKBUF_X2 inst_18556 ( .A(net_18403), .Z(net_18404) );
SDFF_X2 inst_1508 ( .SI(net_7869), .Q(net_7869), .D(net_2660), .SE(net_2558), .CK(net_17011) );
SDFF_X2 inst_1222 ( .Q(net_7956), .D(net_7956), .SE(net_2755), .SI(net_2589), .CK(net_18097) );
AND2_X4 inst_9151 ( .ZN(net_6280), .A2(net_2265), .A1(net_1177) );
CLKBUF_X2 inst_11366 ( .A(net_10602), .Z(net_11214) );
NOR2_X2 inst_3407 ( .ZN(net_3568), .A1(net_3359), .A2(net_3358) );
SDFF_X2 inst_1073 ( .D(net_7321), .SI(net_6497), .Q(net_6497), .SE(net_3071), .CK(net_12092) );
SDFFR_X2 inst_2323 ( .SE(net_2260), .Q(net_376), .D(net_376), .CK(net_9171), .RN(x6501), .SI(x1467) );
NAND4_X2 inst_3741 ( .ZN(net_4289), .A1(net_4070), .A2(net_4069), .A3(net_4068), .A4(net_4067) );
CLKBUF_X2 inst_14643 ( .A(net_14490), .Z(net_14491) );
SDFF_X2 inst_1449 ( .SI(net_7298), .Q(net_7115), .D(net_7115), .SE(net_6278), .CK(net_18200) );
INV_X4 inst_5657 ( .A(net_7354), .ZN(net_1268) );
CLKBUF_X2 inst_11614 ( .A(net_11310), .Z(net_11462) );
AOI22_X2 inst_7872 ( .A2(net_6437), .A1(net_5654), .B2(net_4881), .ZN(net_4569), .B1(net_237) );
XNOR2_X2 inst_187 ( .B(net_6475), .ZN(net_1642), .A(net_1641) );
XNOR2_X2 inst_206 ( .ZN(net_2932), .A(net_2904), .B(net_1508) );
CLKBUF_X2 inst_16449 ( .A(net_16296), .Z(net_16297) );
NAND4_X2 inst_3739 ( .ZN(net_4291), .A1(net_4082), .A2(net_4081), .A3(net_4080), .A4(net_4079) );
SDFF_X2 inst_405 ( .SI(net_8318), .Q(net_8318), .SE(net_3978), .D(net_3956), .CK(net_13291) );
INV_X2 inst_6436 ( .A(net_933), .ZN(net_671) );
NAND2_X2 inst_4788 ( .ZN(net_1532), .A2(net_1136), .A1(net_576) );
CLKBUF_X2 inst_10505 ( .A(net_9347), .Z(net_10353) );
INV_X32 inst_6166 ( .ZN(net_5442), .A(net_4902) );
CLKBUF_X2 inst_17734 ( .A(net_17581), .Z(net_17582) );
CLKBUF_X2 inst_12833 ( .A(net_12680), .Z(net_12681) );
CLKBUF_X2 inst_15868 ( .A(net_15715), .Z(net_15716) );
DFF_X1 inst_6776 ( .Q(net_7555), .D(net_4596), .CK(net_10479) );
CLKBUF_X2 inst_13087 ( .A(net_12934), .Z(net_12935) );
INV_X4 inst_5645 ( .A(net_7207), .ZN(net_1522) );
CLKBUF_X2 inst_18140 ( .A(net_17987), .Z(net_17988) );
CLKBUF_X2 inst_13046 ( .A(net_12893), .Z(net_12894) );
SDFFR_X2 inst_2176 ( .QN(net_7596), .SE(net_3144), .D(net_3113), .SI(net_1011), .CK(net_13495), .RN(x6501) );
OR2_X2 inst_2892 ( .ZN(net_2089), .A1(net_1456), .A2(net_1455) );
INV_X2 inst_6339 ( .A(net_2868), .ZN(net_2691) );
CLKBUF_X2 inst_13024 ( .A(net_12871), .Z(net_12872) );
CLKBUF_X2 inst_19027 ( .A(net_18874), .Z(net_18875) );
CLKBUF_X2 inst_18001 ( .A(net_17848), .Z(net_17849) );
CLKBUF_X2 inst_14929 ( .A(net_12565), .Z(net_14777) );
CLKBUF_X2 inst_15082 ( .A(net_14929), .Z(net_14930) );
CLKBUF_X2 inst_11663 ( .A(net_11510), .Z(net_11511) );
AOI22_X2 inst_7804 ( .A2(net_8221), .B1(net_7177), .B2(net_5655), .A1(net_5268), .ZN(net_4770) );
CLKBUF_X2 inst_14968 ( .A(net_9393), .Z(net_14816) );
CLKBUF_X2 inst_9795 ( .A(net_9642), .Z(net_9643) );
INV_X4 inst_5365 ( .ZN(net_1348), .A(net_1138) );
CLKBUF_X2 inst_15889 ( .A(net_15736), .Z(net_15737) );
SDFFR_X2 inst_2482 ( .Q(net_8988), .D(net_8988), .SI(net_2610), .SE(net_2562), .CK(net_16890), .RN(x6501) );
OAI221_X2 inst_2957 ( .C2(net_8229), .B1(net_7572), .B2(net_4971), .C1(net_4928), .ZN(net_4877), .A(net_3057) );
CLKBUF_X2 inst_15606 ( .A(net_15096), .Z(net_15454) );
CLKBUF_X2 inst_10880 ( .A(net_10523), .Z(net_10728) );
CLKBUF_X2 inst_15551 ( .A(net_15398), .Z(net_15399) );
SDFFR_X1 inst_2711 ( .QN(net_6816), .SE(net_6267), .SI(net_4621), .D(net_1210), .CK(net_11785), .RN(x6501) );
CLKBUF_X2 inst_12808 ( .A(net_12655), .Z(net_12656) );
NOR2_X2 inst_3531 ( .ZN(net_1801), .A2(net_1632), .A1(net_1478) );
SDFFR_X1 inst_2753 ( .QN(net_7573), .D(net_3945), .SE(net_3144), .SI(net_3143), .CK(net_10882), .RN(x6501) );
CLKBUF_X2 inst_16525 ( .A(net_10059), .Z(net_16373) );
NAND4_X2 inst_3672 ( .A4(net_6050), .A1(net_6049), .ZN(net_4593), .A2(net_4060), .A3(net_4059) );
CLKBUF_X2 inst_14329 ( .A(net_14176), .Z(net_14177) );
CLKBUF_X2 inst_16329 ( .A(net_16176), .Z(net_16177) );
XNOR2_X2 inst_132 ( .ZN(net_2815), .B(net_2752), .A(net_2751) );
CLKBUF_X2 inst_18927 ( .A(net_18774), .Z(net_18775) );
CLKBUF_X2 inst_15484 ( .A(net_15331), .Z(net_15332) );
CLKBUF_X2 inst_10353 ( .A(net_10200), .Z(net_10201) );
CLKBUF_X2 inst_13900 ( .A(net_11087), .Z(net_13748) );
CLKBUF_X2 inst_11502 ( .A(net_9751), .Z(net_11350) );
CLKBUF_X2 inst_17092 ( .A(net_16916), .Z(net_16940) );
CLKBUF_X2 inst_12619 ( .A(net_10743), .Z(net_12467) );
CLKBUF_X2 inst_17000 ( .A(net_16847), .Z(net_16848) );
CLKBUF_X2 inst_10369 ( .A(net_10216), .Z(net_10217) );
AOI22_X2 inst_7935 ( .B1(net_7918), .A1(net_7816), .B2(net_6103), .A2(net_4398), .ZN(net_4189) );
INV_X4 inst_6149 ( .A(net_6155), .ZN(net_6154) );
NOR2_X2 inst_3545 ( .A1(net_5974), .ZN(net_1453), .A2(net_1331) );
CLKBUF_X2 inst_16982 ( .A(net_16829), .Z(net_16830) );
CLKBUF_X2 inst_15681 ( .A(net_11544), .Z(net_15529) );
NOR2_X2 inst_3611 ( .A1(net_5967), .A2(net_5966), .ZN(net_2391) );
CLKBUF_X2 inst_12612 ( .A(net_12459), .Z(net_12460) );
CLKBUF_X2 inst_16964 ( .A(net_12916), .Z(net_16812) );
CLKBUF_X2 inst_18476 ( .A(net_18323), .Z(net_18324) );
CLKBUF_X2 inst_17968 ( .A(net_14999), .Z(net_17816) );
CLKBUF_X2 inst_15083 ( .A(net_14431), .Z(net_14931) );
NAND3_X2 inst_3975 ( .ZN(net_2306), .A3(net_1529), .A1(net_796), .A2(net_265) );
CLKBUF_X2 inst_11025 ( .A(net_10394), .Z(net_10873) );
CLKBUF_X2 inst_10976 ( .A(net_10823), .Z(net_10824) );
XNOR2_X2 inst_327 ( .A(net_927), .ZN(net_925), .B(net_196) );
AOI21_X2 inst_8874 ( .ZN(net_5923), .A(net_5922), .B2(net_5843), .B1(x594) );
AOI22_X2 inst_7801 ( .A2(net_6130), .B2(net_4965), .ZN(net_4787), .B1(net_2692), .A1(net_1405) );
CLKBUF_X2 inst_9431 ( .A(net_9278), .Z(net_9279) );
NAND4_X2 inst_3853 ( .ZN(net_1736), .A4(net_1031), .A3(net_977), .A1(net_960), .A2(net_957) );
AOI22_X2 inst_8044 ( .B1(net_8103), .A1(net_7763), .B2(net_6108), .A2(net_6096), .ZN(net_4096) );
CLKBUF_X2 inst_15132 ( .A(net_12878), .Z(net_14980) );
HA_X1 inst_6702 ( .A(net_6220), .CO(net_6078), .S(net_2151), .B(net_2150) );
CLKBUF_X2 inst_14304 ( .A(net_14151), .Z(net_14152) );
CLKBUF_X2 inst_12421 ( .A(net_12268), .Z(net_12269) );
AOI22_X2 inst_7905 ( .B1(net_7192), .A2(net_6443), .B2(net_5655), .A1(net_5654), .ZN(net_4521) );
CLKBUF_X2 inst_17415 ( .A(net_16418), .Z(net_17263) );
CLKBUF_X2 inst_10739 ( .A(net_10586), .Z(net_10587) );
NAND4_X2 inst_3661 ( .A4(net_6040), .A1(net_6039), .ZN(net_4604), .A2(net_4126), .A3(net_4125) );
CLKBUF_X2 inst_16758 ( .A(net_16605), .Z(net_16606) );
CLKBUF_X2 inst_13678 ( .A(net_13525), .Z(net_13526) );
CLKBUF_X2 inst_14244 ( .A(net_14091), .Z(net_14092) );
CLKBUF_X2 inst_15963 ( .A(net_14190), .Z(net_15811) );
AOI21_X2 inst_9001 ( .B1(net_7353), .ZN(net_1270), .A(net_1269), .B2(net_1268) );
CLKBUF_X2 inst_11836 ( .A(net_9938), .Z(net_11684) );
NOR4_X2 inst_3221 ( .ZN(net_2491), .A3(net_2295), .A4(net_2291), .A1(net_1299), .A2(net_1297) );
CLKBUF_X2 inst_16251 ( .A(net_16098), .Z(net_16099) );
CLKBUF_X2 inst_14585 ( .A(net_13340), .Z(net_14433) );
CLKBUF_X2 inst_16209 ( .A(net_11989), .Z(net_16057) );
CLKBUF_X2 inst_12335 ( .A(net_9763), .Z(net_12183) );
SDFF_X2 inst_357 ( .Q(net_8760), .D(net_8760), .SE(net_3982), .SI(net_3974), .CK(net_10863) );
CLKBUF_X2 inst_11083 ( .A(net_10930), .Z(net_10931) );
DFFR_X2 inst_6969 ( .QN(net_5971), .D(net_5926), .CK(net_11566), .RN(x6501) );
CLKBUF_X2 inst_10028 ( .A(net_9875), .Z(net_9876) );
INV_X2 inst_6173 ( .ZN(net_5932), .A(net_5924) );
NAND2_X2 inst_4092 ( .ZN(net_5446), .A1(net_5167), .A2(net_5165) );
CLKBUF_X2 inst_13865 ( .A(net_13712), .Z(net_13713) );
CLKBUF_X2 inst_10098 ( .A(net_9945), .Z(net_9946) );
NAND3_X2 inst_3980 ( .ZN(net_2387), .A3(net_2315), .A2(net_1881), .A1(net_1781) );
CLKBUF_X2 inst_11438 ( .A(net_9305), .Z(net_11286) );
NAND4_X2 inst_3758 ( .A3(net_6075), .A1(net_6074), .ZN(net_4263), .A2(net_3842), .A4(net_3841) );
SDFF_X2 inst_912 ( .SI(net_8731), .Q(net_8731), .SE(net_6195), .D(net_3941), .CK(net_10316) );
CLKBUF_X2 inst_18087 ( .A(net_17934), .Z(net_17935) );
CLKBUF_X2 inst_15653 ( .A(net_15500), .Z(net_15501) );
CLKBUF_X2 inst_10065 ( .A(net_9912), .Z(net_9913) );
CLKBUF_X2 inst_15923 ( .A(net_9969), .Z(net_15771) );
CLKBUF_X2 inst_18516 ( .A(net_18363), .Z(net_18364) );
CLKBUF_X2 inst_18451 ( .A(net_16548), .Z(net_18299) );
CLKBUF_X2 inst_12724 ( .A(net_12571), .Z(net_12572) );
INV_X4 inst_5872 ( .A(net_8938), .ZN(net_4743) );
CLKBUF_X2 inst_16735 ( .A(net_16582), .Z(net_16583) );
DFFR_X2 inst_6988 ( .QN(net_5961), .D(net_5899), .CK(net_11493), .RN(x6501) );
NAND2_X2 inst_4188 ( .ZN(net_5313), .A1(net_5068), .A2(net_5067) );
CLKBUF_X2 inst_14888 ( .A(net_14735), .Z(net_14736) );
CLKBUF_X2 inst_14405 ( .A(net_9970), .Z(net_14253) );
NAND2_X2 inst_4169 ( .ZN(net_5341), .A1(net_5197), .A2(net_4991) );
CLKBUF_X2 inst_16755 ( .A(net_16602), .Z(net_16603) );
CLKBUF_X2 inst_9894 ( .A(net_9306), .Z(net_9742) );
DFFS_X2 inst_6863 ( .Q(net_6322), .D(net_5532), .CK(net_18935), .SN(x6501) );
CLKBUF_X2 inst_18149 ( .A(net_17996), .Z(net_17997) );
INV_X4 inst_5346 ( .ZN(net_2008), .A(net_1910) );
NAND2_X2 inst_4181 ( .ZN(net_5322), .A1(net_5189), .A2(net_4987) );
CLKBUF_X2 inst_10865 ( .A(net_10340), .Z(net_10713) );
SDFF_X2 inst_2008 ( .SI(net_7796), .Q(net_7796), .D(net_2717), .SE(net_2459), .CK(net_16456) );
CLKBUF_X2 inst_16786 ( .A(net_16633), .Z(net_16634) );
SDFF_X2 inst_641 ( .SI(net_8523), .Q(net_8523), .SE(net_3979), .D(net_3938), .CK(net_12974) );
SDFF_X2 inst_498 ( .SI(net_8623), .Q(net_8623), .SE(net_3984), .D(net_3940), .CK(net_13483) );
CLKBUF_X2 inst_17902 ( .A(net_17749), .Z(net_17750) );
CLKBUF_X2 inst_17623 ( .A(net_17470), .Z(net_17471) );
SDFF_X2 inst_1988 ( .D(net_7282), .SI(net_7019), .Q(net_7019), .SE(net_6277), .CK(net_14867) );
AOI22_X2 inst_8374 ( .B1(net_8855), .A1(net_8300), .B2(net_6252), .A2(net_4345), .ZN(net_3674) );
CLKBUF_X2 inst_12346 ( .A(net_12193), .Z(net_12194) );
AOI22_X2 inst_8287 ( .B1(net_8730), .A1(net_8508), .B2(net_4350), .A2(net_4349), .ZN(net_3755) );
CLKBUF_X2 inst_11971 ( .A(net_11628), .Z(net_11819) );
INV_X4 inst_5517 ( .ZN(net_880), .A(net_676) );
SDFF_X2 inst_1912 ( .D(net_7286), .SI(net_6863), .Q(net_6863), .SE(net_6282), .CK(net_16174) );
CLKBUF_X2 inst_14478 ( .A(net_13920), .Z(net_14326) );
SDFF_X2 inst_1831 ( .D(net_7295), .SI(net_6872), .Q(net_6872), .SE(net_6282), .CK(net_15416) );
CLKBUF_X2 inst_13438 ( .A(net_13285), .Z(net_13286) );
HA_X1 inst_6714 ( .A(net_3600), .B(net_3595), .CO(net_1567), .S(net_1229) );
HA_X1 inst_6683 ( .S(net_3016), .CO(net_3015), .A(net_3014), .B(net_2819) );
CLKBUF_X2 inst_14339 ( .A(net_12712), .Z(net_14187) );
CLKBUF_X2 inst_13671 ( .A(net_13518), .Z(net_13519) );
NOR2_X2 inst_3468 ( .ZN(net_2554), .A2(net_2464), .A1(net_2457) );
SDFFR_X2 inst_2395 ( .SE(net_2260), .Q(net_351), .D(net_351), .CK(net_9287), .RN(x6501), .SI(x2230) );
XNOR2_X2 inst_231 ( .ZN(net_1299), .A(net_1298), .B(net_776) );
AND4_X4 inst_9024 ( .ZN(net_4970), .A4(net_4722), .A1(net_4581), .A2(net_4546), .A3(net_4483) );
NOR3_X2 inst_3309 ( .ZN(net_1742), .A1(net_1224), .A2(net_1088), .A3(net_1010) );
CLKBUF_X2 inst_9952 ( .A(net_9799), .Z(net_9800) );
INV_X4 inst_5676 ( .A(net_6394), .ZN(net_2141) );
CLKBUF_X2 inst_15459 ( .A(net_12450), .Z(net_15307) );
SDFFR_X2 inst_2317 ( .QN(net_7477), .SE(net_3354), .SI(net_3129), .CK(net_9970), .D(x13364), .RN(x6501) );
CLKBUF_X2 inst_11365 ( .A(net_11212), .Z(net_11213) );
CLKBUF_X2 inst_15816 ( .A(net_15663), .Z(net_15664) );
DFF_X1 inst_6756 ( .Q(net_7527), .D(net_4616), .CK(net_9543) );
CLKBUF_X2 inst_15208 ( .A(net_10420), .Z(net_15056) );
MUX2_X2 inst_5000 ( .A(net_9039), .Z(net_3955), .B(net_3227), .S(net_622) );
NAND2_X2 inst_4077 ( .A2(net_6779), .A1(net_5835), .ZN(net_5769) );
OAI21_X2 inst_3139 ( .B2(net_2060), .ZN(net_2058), .A(net_1968), .B1(net_606) );
CLKBUF_X2 inst_12801 ( .A(net_9709), .Z(net_12649) );
SDFFR_X2 inst_2558 ( .SI(net_7262), .Q(net_6383), .D(net_6383), .SE(net_2147), .CK(net_15032), .RN(x6501) );
CLKBUF_X2 inst_18591 ( .A(net_14807), .Z(net_18439) );
SDFF_X2 inst_352 ( .SI(net_8455), .Q(net_8455), .SE(net_3983), .D(net_3960), .CK(net_13379) );
XNOR2_X2 inst_286 ( .A(net_1776), .ZN(net_1009), .B(net_199) );
CLKBUF_X2 inst_17452 ( .A(net_17299), .Z(net_17300) );
CLKBUF_X2 inst_13354 ( .A(net_9901), .Z(net_13202) );
CLKBUF_X2 inst_10112 ( .A(net_9959), .Z(net_9960) );
DFFS_X2 inst_6880 ( .Q(net_6324), .D(net_3214), .CK(net_14473), .SN(x6501) );
CLKBUF_X2 inst_15328 ( .A(net_15175), .Z(net_15176) );
CLKBUF_X2 inst_15663 ( .A(net_15510), .Z(net_15511) );
CLKBUF_X2 inst_10447 ( .A(net_10294), .Z(net_10295) );
CLKBUF_X2 inst_14959 ( .A(net_14806), .Z(net_14807) );
CLKBUF_X2 inst_12984 ( .A(net_12831), .Z(net_12832) );
CLKBUF_X2 inst_15524 ( .A(net_15371), .Z(net_15372) );
CLKBUF_X2 inst_13006 ( .A(net_12853), .Z(net_12854) );
AOI22_X2 inst_7961 ( .B1(net_8126), .A1(net_7888), .A2(net_6098), .B2(net_4190), .ZN(net_4167) );
CLKBUF_X2 inst_16900 ( .A(net_16747), .Z(net_16748) );
DFF_X1 inst_6792 ( .Q(net_8239), .D(net_4441), .CK(net_14467) );
CLKBUF_X2 inst_16361 ( .A(net_11720), .Z(net_16209) );
CLKBUF_X2 inst_15058 ( .A(net_14905), .Z(net_14906) );
NAND4_X2 inst_3841 ( .ZN(net_2112), .A2(net_1654), .A1(net_1172), .A4(net_151), .A3(net_150) );
CLKBUF_X2 inst_9555 ( .A(net_9223), .Z(net_9403) );
AOI22_X4 inst_7737 ( .A2(net_8613), .B1(net_8428), .A1(net_3864), .B2(net_3863), .ZN(net_3787) );
DFFR_X2 inst_6972 ( .QN(net_7622), .D(net_5929), .CK(net_11180), .RN(x6501) );
CLKBUF_X2 inst_12203 ( .A(net_12050), .Z(net_12051) );
CLKBUF_X2 inst_9427 ( .A(net_9274), .Z(net_9275) );
INV_X4 inst_5887 ( .A(net_6836), .ZN(net_681) );
CLKBUF_X2 inst_11598 ( .A(net_10093), .Z(net_11446) );
CLKBUF_X2 inst_13452 ( .A(net_13299), .Z(net_13300) );
CLKBUF_X2 inst_12001 ( .A(net_11848), .Z(net_11849) );
CLKBUF_X2 inst_17809 ( .A(net_17656), .Z(net_17657) );
SDFF_X2 inst_425 ( .Q(net_8751), .D(net_8751), .SE(net_3982), .SI(net_3960), .CK(net_13151) );
AOI22_X2 inst_8416 ( .B1(net_8861), .A1(net_8306), .B2(net_6252), .A2(net_4345), .ZN(net_3636) );
CLKBUF_X2 inst_15298 ( .A(net_15145), .Z(net_15146) );
SDFFR_X2 inst_2572 ( .QN(net_6350), .SE(net_2147), .D(net_2079), .SI(net_1854), .CK(net_17519), .RN(x6501) );
CLKBUF_X2 inst_13764 ( .A(net_11357), .Z(net_13612) );
CLKBUF_X2 inst_9380 ( .A(net_9227), .Z(net_9228) );
DFF_X1 inst_6755 ( .Q(net_7645), .D(net_4590), .CK(net_10801) );
CLKBUF_X2 inst_13111 ( .A(net_12958), .Z(net_12959) );
NOR2_X2 inst_3365 ( .ZN(net_5560), .A1(net_5368), .A2(net_5367) );
NOR3_X2 inst_3254 ( .ZN(net_5453), .A1(net_5452), .A3(net_4938), .A2(net_2900) );
CLKBUF_X2 inst_17885 ( .A(net_17732), .Z(net_17733) );
SDFF_X2 inst_983 ( .SI(net_7320), .Q(net_6727), .D(net_6727), .SE(net_3124), .CK(net_9876) );
MUX2_X2 inst_4980 ( .A(net_9044), .B(net_7441), .Z(net_3952), .S(net_622) );
AOI22_X2 inst_8026 ( .B1(net_7930), .A1(net_7828), .B2(net_6103), .A2(net_4398), .ZN(net_4111) );
AOI22_X2 inst_7773 ( .B1(net_6963), .A1(net_6923), .A2(net_5443), .B2(net_5442), .ZN(net_5311) );
CLKBUF_X2 inst_17426 ( .A(net_17273), .Z(net_17274) );
CLKBUF_X2 inst_11291 ( .A(net_11138), .Z(net_11139) );
CLKBUF_X2 inst_11196 ( .A(net_11043), .Z(net_11044) );
NAND2_X2 inst_4776 ( .A2(net_7220), .ZN(net_1803), .A1(net_1631) );
INV_X2 inst_6237 ( .ZN(net_5282), .A(net_5035) );
SDFFR_X2 inst_2633 ( .Q(net_7383), .D(net_7383), .SE(net_1136), .CK(net_18608), .RN(x6501), .SI(x4693) );
DFFS_X1 inst_6947 ( .D(net_6145), .CK(net_13630), .SN(x6501), .Q(x735) );
INV_X2 inst_6274 ( .ZN(net_4377), .A(net_4363) );
DFFR_X2 inst_7029 ( .QN(net_7208), .D(net_5592), .CK(net_18965), .RN(x6501) );
SDFFR_X2 inst_2130 ( .SI(net_7195), .Q(net_7195), .D(net_6446), .SE(net_4362), .CK(net_13561), .RN(x6501) );
NAND2_X2 inst_4388 ( .A1(net_7079), .A2(net_5162), .ZN(net_5069) );
SDFF_X2 inst_1055 ( .SI(net_7323), .Q(net_6664), .D(net_6664), .SE(net_3126), .CK(net_9133) );
CLKBUF_X2 inst_13114 ( .A(net_9215), .Z(net_12962) );
SDFFS_X1 inst_2100 ( .SI(net_6817), .Q(net_6817), .SE(net_6269), .D(net_1208), .CK(net_11775), .SN(x6501) );
CLKBUF_X2 inst_16813 ( .A(net_14865), .Z(net_16661) );
SDFFR_X2 inst_2284 ( .SE(net_2789), .SI(net_2760), .Q(net_256), .D(net_256), .CK(net_13706), .RN(x6501) );
CLKBUF_X2 inst_16028 ( .A(net_15875), .Z(net_15876) );
NAND2_X2 inst_4829 ( .A1(net_4890), .ZN(net_1320), .A2(net_1099) );
CLKBUF_X2 inst_16032 ( .A(net_15267), .Z(net_15880) );
CLKBUF_X2 inst_16505 ( .A(net_14021), .Z(net_16353) );
CLKBUF_X2 inst_19041 ( .A(net_18888), .Z(net_18889) );
SDFF_X2 inst_923 ( .SI(net_8711), .Q(net_8711), .SE(net_6195), .D(net_3981), .CK(net_12940) );
CLKBUF_X2 inst_12153 ( .A(net_12000), .Z(net_12001) );
AOI222_X1 inst_8671 ( .C2(net_5832), .A2(net_5830), .B2(net_5824), .ZN(net_3584), .A1(net_3279), .B1(net_2144), .C1(x2355) );
AOI222_X1 inst_8599 ( .B2(net_6781), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5826), .A1(net_3580), .C1(x2494) );
CLKBUF_X2 inst_17569 ( .A(net_17416), .Z(net_17417) );
CLKBUF_X2 inst_11604 ( .A(net_11451), .Z(net_11452) );
CLKBUF_X2 inst_13470 ( .A(net_13317), .Z(net_13318) );
DFFR_X2 inst_6975 ( .QN(net_5963), .D(net_5909), .CK(net_9348), .RN(x6501) );
CLKBUF_X2 inst_11819 ( .A(net_9211), .Z(net_11667) );
DFFR_X1 inst_7564 ( .D(net_7667), .Q(net_7655), .CK(net_12699), .RN(x6501) );
DFFR_X2 inst_7109 ( .QN(net_7635), .D(net_3155), .CK(net_18957), .RN(x6501) );
CLKBUF_X2 inst_16073 ( .A(net_15920), .Z(net_15921) );
INV_X4 inst_5890 ( .A(net_5960), .ZN(x2856) );
CLKBUF_X2 inst_18764 ( .A(net_18611), .Z(net_18612) );
AOI221_X2 inst_8793 ( .B1(net_5268), .ZN(net_4906), .A(net_4905), .B2(net_4627), .C2(net_4388), .C1(net_2614) );
CLKBUF_X2 inst_12946 ( .A(net_12793), .Z(net_12794) );
NAND4_X2 inst_3766 ( .ZN(net_4255), .A1(net_3790), .A2(net_3789), .A3(net_3788), .A4(net_3787) );
CLKBUF_X2 inst_12480 ( .A(net_12300), .Z(net_12328) );
INV_X4 inst_5935 ( .A(net_7236), .ZN(net_1866) );
SDFFR_X2 inst_2536 ( .QN(net_6353), .SE(net_2147), .D(net_2145), .SI(net_1855), .CK(net_17537), .RN(x6501) );
CLKBUF_X2 inst_11730 ( .A(net_11577), .Z(net_11578) );
CLKBUF_X2 inst_13103 ( .A(net_12766), .Z(net_12951) );
CLKBUF_X2 inst_9389 ( .A(net_9236), .Z(net_9237) );
DFFR_X2 inst_7100 ( .QN(net_5978), .D(net_3261), .CK(net_11232), .RN(x6501) );
CLKBUF_X2 inst_9618 ( .A(net_9465), .Z(net_9466) );
CLKBUF_X2 inst_14036 ( .A(net_12569), .Z(net_13884) );
DFFS_X2 inst_6870 ( .QN(net_8293), .D(net_4224), .CK(net_11207), .SN(x6501) );
CLKBUF_X2 inst_13300 ( .A(net_9303), .Z(net_13148) );
INV_X4 inst_5915 ( .A(net_7502), .ZN(net_3272) );
CLKBUF_X2 inst_10998 ( .A(net_10845), .Z(net_10846) );
SDFF_X2 inst_1925 ( .D(net_7264), .SI(net_6881), .Q(net_6881), .SE(net_6284), .CK(net_14323) );
XOR2_X2 inst_40 ( .A(net_3048), .Z(net_1048), .B(net_536) );
NAND2_X2 inst_4437 ( .A1(net_6874), .A2(net_5016), .ZN(net_4990) );
CLKBUF_X2 inst_16007 ( .A(net_15854), .Z(net_15855) );
AOI221_X2 inst_8765 ( .C2(net_5657), .B2(net_5463), .ZN(net_5460), .A(net_4942), .C1(net_2700), .B1(net_434) );
SDFF_X2 inst_1416 ( .SI(net_7296), .Q(net_7153), .D(net_7153), .SE(net_6279), .CK(net_18211) );
CLKBUF_X2 inst_12066 ( .A(net_10212), .Z(net_11914) );
DFFR_X2 inst_7280 ( .QN(net_6390), .D(net_1768), .CK(net_15662), .RN(x6501) );
SDFF_X2 inst_439 ( .Q(net_8768), .D(net_8768), .SE(net_3982), .SI(net_3941), .CK(net_10383) );
CLKBUF_X2 inst_17304 ( .A(net_15138), .Z(net_17152) );
CLKBUF_X2 inst_16582 ( .A(net_16429), .Z(net_16430) );
CLKBUF_X2 inst_11567 ( .A(net_11414), .Z(net_11415) );
NAND2_X2 inst_4529 ( .A2(net_3574), .ZN(net_3556), .A1(net_3555) );
CLKBUF_X2 inst_17445 ( .A(net_17292), .Z(net_17293) );
CLKBUF_X2 inst_15216 ( .A(net_15063), .Z(net_15064) );
AOI22_X2 inst_8280 ( .B1(net_8803), .A1(net_8544), .A2(net_3861), .B2(net_3860), .ZN(net_3761) );
CLKBUF_X2 inst_16816 ( .A(net_16663), .Z(net_16664) );
CLKBUF_X2 inst_13309 ( .A(net_13156), .Z(net_13157) );
CLKBUF_X2 inst_13475 ( .A(net_13322), .Z(net_13323) );
CLKBUF_X2 inst_17009 ( .A(net_10550), .Z(net_16857) );
CLKBUF_X2 inst_9478 ( .A(net_9325), .Z(net_9326) );
CLKBUF_X2 inst_18643 ( .A(net_18490), .Z(net_18491) );
SDFF_X2 inst_654 ( .Q(net_8427), .D(net_8427), .SI(net_3974), .SE(net_3934), .CK(net_10830) );
CLKBUF_X2 inst_17077 ( .A(net_12892), .Z(net_16925) );
CLKBUF_X2 inst_16152 ( .A(net_12399), .Z(net_16000) );
CLKBUF_X2 inst_13616 ( .A(net_12521), .Z(net_13464) );
CLKBUF_X2 inst_16284 ( .A(net_16131), .Z(net_16132) );
CLKBUF_X2 inst_16486 ( .A(net_16333), .Z(net_16334) );
CLKBUF_X2 inst_13656 ( .A(net_12258), .Z(net_13504) );
CLKBUF_X2 inst_17130 ( .A(net_16977), .Z(net_16978) );
CLKBUF_X2 inst_16574 ( .A(net_16421), .Z(net_16422) );
SDFF_X2 inst_1708 ( .Q(net_8009), .D(net_8009), .SI(net_2703), .SE(net_2542), .CK(net_16713) );
CLKBUF_X2 inst_15264 ( .A(net_9699), .Z(net_15112) );
CLKBUF_X2 inst_15096 ( .A(net_12139), .Z(net_14944) );
CLKBUF_X2 inst_11997 ( .A(net_9743), .Z(net_11845) );
CLKBUF_X2 inst_10440 ( .A(net_9763), .Z(net_10288) );
CLKBUF_X2 inst_11004 ( .A(net_10851), .Z(net_10852) );
CLKBUF_X2 inst_17469 ( .A(net_17316), .Z(net_17317) );
SDFFR_X1 inst_2738 ( .SI(net_9020), .Q(net_9020), .D(net_7449), .SE(net_3208), .CK(net_10101), .RN(x6501) );
CLKBUF_X2 inst_16164 ( .A(net_15455), .Z(net_16012) );
SDFF_X2 inst_634 ( .SI(net_8548), .Q(net_8548), .SE(net_3979), .D(net_3952), .CK(net_12884) );
OAI21_X2 inst_3122 ( .B1(net_6837), .ZN(net_2285), .A(net_2283), .B2(net_2282) );
CLKBUF_X2 inst_15229 ( .A(net_15076), .Z(net_15077) );
AND2_X4 inst_9090 ( .A2(net_2440), .ZN(net_2439), .A1(net_2342) );
CLKBUF_X2 inst_16989 ( .A(net_16836), .Z(net_16837) );
CLKBUF_X2 inst_17184 ( .A(net_17031), .Z(net_17032) );
CLKBUF_X2 inst_9232 ( .A(net_9079), .Z(net_9080) );
CLKBUF_X2 inst_10420 ( .A(net_10267), .Z(net_10268) );
CLKBUF_X2 inst_18202 ( .A(net_18049), .Z(net_18050) );
SDFF_X2 inst_1477 ( .SI(net_7272), .Q(net_7129), .D(net_7129), .SE(net_6279), .CK(net_16837) );
CLKBUF_X2 inst_13774 ( .A(net_9523), .Z(net_13622) );
CLKBUF_X2 inst_9263 ( .A(net_9110), .Z(net_9111) );
DFFR_X2 inst_7043 ( .QN(net_7501), .D(net_4929), .CK(net_16681), .RN(x6501) );
CLKBUF_X2 inst_9813 ( .A(net_9660), .Z(net_9661) );
SDFF_X2 inst_529 ( .Q(net_8885), .D(net_8885), .SI(net_3976), .SE(net_3936), .CK(net_12897) );
SDFF_X2 inst_1528 ( .Q(net_7904), .D(net_7904), .SI(net_2704), .SE(net_2543), .CK(net_14279) );
CLKBUF_X2 inst_11192 ( .A(net_11039), .Z(net_11040) );
CLKBUF_X2 inst_17122 ( .A(net_16969), .Z(net_16970) );
CLKBUF_X2 inst_15921 ( .A(net_9292), .Z(net_15769) );
CLKBUF_X2 inst_15705 ( .A(net_15552), .Z(net_15553) );
CLKBUF_X2 inst_16333 ( .A(net_16180), .Z(net_16181) );
INV_X4 inst_5788 ( .A(net_7521), .ZN(net_1076) );
CLKBUF_X2 inst_11788 ( .A(net_9929), .Z(net_11636) );
CLKBUF_X2 inst_17562 ( .A(net_9135), .Z(net_17410) );
CLKBUF_X2 inst_15460 ( .A(net_15307), .Z(net_15308) );
CLKBUF_X2 inst_14267 ( .A(net_12126), .Z(net_14115) );
CLKBUF_X2 inst_11030 ( .A(net_9079), .Z(net_10878) );
SDFF_X2 inst_675 ( .Q(net_8673), .D(net_8673), .SI(net_3947), .SE(net_3935), .CK(net_12963) );
NAND2_X2 inst_4068 ( .ZN(net_5840), .A2(net_5764), .A1(net_3210) );
CLKBUF_X2 inst_11953 ( .A(net_11800), .Z(net_11801) );
CLKBUF_X2 inst_13706 ( .A(net_9554), .Z(net_13554) );
INV_X4 inst_5729 ( .A(net_8931), .ZN(net_2604) );
SDFFR_X1 inst_2705 ( .SI(net_6814), .Q(net_6814), .D(net_6811), .SE(net_6268), .CK(net_11799), .RN(x6501) );
CLKBUF_X2 inst_19192 ( .A(net_19039), .Z(net_19040) );
CLKBUF_X2 inst_16662 ( .A(net_16509), .Z(net_16510) );
CLKBUF_X2 inst_13291 ( .A(net_13138), .Z(net_13139) );
CLKBUF_X2 inst_12902 ( .A(net_12749), .Z(net_12750) );
CLKBUF_X2 inst_12924 ( .A(net_12771), .Z(net_12772) );
INV_X4 inst_5737 ( .A(net_6300), .ZN(net_2689) );
INV_X4 inst_5332 ( .ZN(net_1477), .A(net_1344) );
CLKBUF_X2 inst_11144 ( .A(net_10194), .Z(net_10992) );
AND2_X4 inst_9078 ( .A2(net_6198), .ZN(net_5830), .A1(net_2986) );
NAND4_X2 inst_3751 ( .ZN(net_4279), .A1(net_4008), .A2(net_4007), .A3(net_4006), .A4(net_4005) );
CLKBUF_X2 inst_17272 ( .A(net_17119), .Z(net_17120) );
CLKBUF_X2 inst_12463 ( .A(net_10358), .Z(net_12311) );
DFF_X1 inst_6735 ( .Q(net_6780), .D(net_5634), .CK(net_9204) );
INV_X16 inst_6643 ( .ZN(net_3867), .A(net_3313) );
CLKBUF_X2 inst_16538 ( .A(net_16385), .Z(net_16386) );
AND2_X4 inst_9123 ( .A1(net_7216), .ZN(net_1836), .A2(net_1089) );
SDFFR_X2 inst_2222 ( .Q(net_7450), .D(net_7450), .SE(net_2863), .CK(net_12812), .SI(x13576), .RN(x6501) );
NAND2_X2 inst_4578 ( .ZN(net_2960), .A1(net_2959), .A2(net_2952) );
CLKBUF_X2 inst_12102 ( .A(net_11949), .Z(net_11950) );
NAND2_X2 inst_4059 ( .ZN(net_5882), .A2(net_5771), .A1(net_3202) );
SDFF_X2 inst_1755 ( .SI(net_7288), .Q(net_7145), .D(net_7145), .SE(net_6279), .CK(net_14903) );
CLKBUF_X2 inst_15390 ( .A(net_15237), .Z(net_15238) );
CLKBUF_X2 inst_15027 ( .A(net_12081), .Z(net_14875) );
CLKBUF_X2 inst_12715 ( .A(net_12562), .Z(net_12563) );
SDFF_X2 inst_806 ( .SI(net_8495), .Q(net_8495), .D(net_3966), .SE(net_3884), .CK(net_9984) );
CLKBUF_X2 inst_18851 ( .A(net_18698), .Z(net_18699) );
DFFR_X2 inst_7119 ( .Q(net_7616), .D(net_3095), .CK(net_11165), .RN(x6501) );
DFFR_X2 inst_7232 ( .QN(net_8216), .D(net_2176), .CK(net_17305), .RN(x6501) );
SDFF_X2 inst_491 ( .SI(net_8615), .Q(net_8615), .SE(net_3984), .D(net_3963), .CK(net_10941) );
CLKBUF_X2 inst_10485 ( .A(net_9154), .Z(net_10333) );
INV_X4 inst_6027 ( .A(net_7513), .ZN(net_506) );
MUX2_X2 inst_4943 ( .B(net_6319), .S(net_5522), .Z(net_2636), .A(net_2635) );
CLKBUF_X2 inst_13219 ( .A(net_13066), .Z(net_13067) );
CLKBUF_X2 inst_13515 ( .A(net_13362), .Z(net_13363) );
CLKBUF_X2 inst_10987 ( .A(net_10834), .Z(net_10835) );
CLKBUF_X2 inst_12097 ( .A(net_11944), .Z(net_11945) );
CLKBUF_X2 inst_9441 ( .A(net_9264), .Z(net_9289) );
OAI21_X2 inst_3086 ( .ZN(net_3157), .B2(net_3033), .A(net_2950), .B1(net_516) );
SDFFR_X1 inst_2791 ( .Q(net_7294), .D(net_2760), .SI(net_1947), .SE(net_1327), .CK(net_15356), .RN(x6501) );
CLKBUF_X2 inst_12090 ( .A(net_11937), .Z(net_11938) );
INV_X4 inst_5583 ( .A(net_7161), .ZN(net_635) );
CLKBUF_X2 inst_16514 ( .A(net_9513), .Z(net_16362) );
CLKBUF_X2 inst_10243 ( .A(net_9758), .Z(net_10091) );
CLKBUF_X2 inst_15633 ( .A(net_15480), .Z(net_15481) );
CLKBUF_X2 inst_14814 ( .A(net_14661), .Z(net_14662) );
NAND2_X2 inst_4419 ( .A1(net_6858), .A2(net_5016), .ZN(net_5008) );
CLKBUF_X2 inst_16342 ( .A(net_16189), .Z(net_16190) );
DFF_X1 inst_6850 ( .Q(net_6438), .D(net_3631), .CK(net_17898) );
HA_X1 inst_6698 ( .S(net_2566), .CO(net_2565), .B(net_2504), .A(x3156) );
SDFF_X2 inst_1349 ( .SI(net_7754), .Q(net_7754), .D(net_2575), .SE(net_2560), .CK(net_16004) );
CLKBUF_X2 inst_18390 ( .A(net_18237), .Z(net_18238) );
DFFR_X2 inst_7012 ( .QN(net_9012), .D(net_5782), .CK(net_11175), .RN(x6501) );
CLKBUF_X2 inst_12744 ( .A(net_12591), .Z(net_12592) );
NAND4_X2 inst_3745 ( .ZN(net_4285), .A1(net_4046), .A2(net_4045), .A3(net_4044), .A4(net_4043) );
CLKBUF_X2 inst_15345 ( .A(net_15192), .Z(net_15193) );
NAND2_X2 inst_4347 ( .A1(net_7147), .A2(net_5166), .ZN(net_5110) );
CLKBUF_X2 inst_16404 ( .A(net_9062), .Z(net_16252) );
INV_X4 inst_5962 ( .A(net_7439), .ZN(net_3533) );
SDFFR_X2 inst_2224 ( .Q(net_7475), .D(net_7475), .SE(net_2863), .CK(net_12186), .SI(x13385), .RN(x6501) );
CLKBUF_X2 inst_10002 ( .A(net_9849), .Z(net_9850) );
CLKBUF_X2 inst_10185 ( .A(net_10032), .Z(net_10033) );
INV_X4 inst_5226 ( .ZN(net_2275), .A(net_2201) );
CLKBUF_X2 inst_13012 ( .A(net_12859), .Z(net_12860) );
INV_X4 inst_5310 ( .A(net_1507), .ZN(net_1476) );
AOI22_X2 inst_8412 ( .B1(net_8750), .A1(net_8380), .A2(net_3867), .B2(net_3866), .ZN(net_3640) );
MUX2_X2 inst_4996 ( .A(net_9030), .Z(net_3973), .B(net_3048), .S(net_622) );
SDFF_X2 inst_1890 ( .D(net_7273), .SI(net_7010), .Q(net_7010), .SE(net_6277), .CK(net_14098) );
SDFFR_X2 inst_2308 ( .SI(net_7406), .SE(net_2260), .Q(net_343), .D(net_343), .CK(net_9369), .RN(x6501) );
NAND2_X2 inst_4093 ( .ZN(net_5445), .A2(net_5250), .A1(net_5163) );
OR2_X2 inst_2879 ( .ZN(net_3063), .A2(net_2881), .A1(net_2835) );
CLKBUF_X2 inst_14676 ( .A(net_14523), .Z(net_14524) );
DFFR_X1 inst_7482 ( .QN(net_7434), .D(net_4210), .CK(net_10113), .RN(x6501) );
SDFFR_X2 inst_2338 ( .SE(net_2260), .Q(net_362), .D(net_362), .CK(net_9315), .RN(x6501), .SI(x1885) );
NOR2_X2 inst_3475 ( .ZN(net_2480), .A2(net_2198), .A1(net_1098) );
CLKBUF_X2 inst_13170 ( .A(net_13017), .Z(net_13018) );
CLKBUF_X2 inst_15547 ( .A(net_15394), .Z(net_15395) );
AOI22_X2 inst_7818 ( .A2(net_8219), .A1(net_5268), .ZN(net_4733), .B1(net_4732), .B2(net_4388) );
CLKBUF_X2 inst_11431 ( .A(net_10630), .Z(net_11279) );
CLKBUF_X2 inst_18319 ( .A(net_18166), .Z(net_18167) );
CLKBUF_X2 inst_18977 ( .A(net_18824), .Z(net_18825) );
INV_X2 inst_6516 ( .ZN(net_889), .A(net_208) );
AOI222_X1 inst_8649 ( .A2(net_6266), .C2(net_6215), .C1(net_4365), .B2(net_4364), .ZN(net_3917), .B1(net_1039), .A1(x13969) );
INV_X4 inst_5198 ( .ZN(net_2495), .A(net_2456) );
INV_X4 inst_5909 ( .A(net_6799), .ZN(net_4360) );
CLKBUF_X2 inst_19003 ( .A(net_16658), .Z(net_18851) );
CLKBUF_X2 inst_16341 ( .A(net_16188), .Z(net_16189) );
CLKBUF_X2 inst_15934 ( .A(net_15781), .Z(net_15782) );
SDFF_X2 inst_2016 ( .SI(net_7794), .Q(net_7794), .D(net_2712), .SE(net_2459), .CK(net_14239) );
CLKBUF_X2 inst_15679 ( .A(net_15526), .Z(net_15527) );
CLKBUF_X2 inst_12723 ( .A(net_12570), .Z(net_12571) );
CLKBUF_X2 inst_16431 ( .A(net_16278), .Z(net_16279) );
NAND3_X1 inst_4012 ( .ZN(net_1306), .A3(x13263), .A1(x13252), .A2(x13234) );
AOI22_X2 inst_8385 ( .B1(net_8783), .A1(net_8524), .A2(net_3861), .B2(net_3860), .ZN(net_3663) );
CLKBUF_X2 inst_15152 ( .A(net_14999), .Z(net_15000) );
CLKBUF_X2 inst_9289 ( .A(net_9136), .Z(net_9137) );
CLKBUF_X2 inst_9920 ( .A(net_9767), .Z(net_9768) );
SDFF_X2 inst_393 ( .Q(net_8834), .D(net_8834), .SI(net_3974), .SE(net_3964), .CK(net_10854) );
INV_X4 inst_5969 ( .A(net_7575), .ZN(net_514) );
SDFF_X2 inst_1813 ( .D(net_7301), .SI(net_6878), .Q(net_6878), .SE(net_6282), .CK(net_15879) );
XOR2_X1 inst_92 ( .Z(net_1418), .B(net_1417), .A(net_651) );
CLKBUF_X2 inst_15405 ( .A(net_15252), .Z(net_15253) );
CLKBUF_X2 inst_11168 ( .A(net_9265), .Z(net_11016) );
SDFF_X2 inst_345 ( .SI(net_8477), .Q(net_8477), .SE(net_3983), .D(net_3950), .CK(net_11030) );
CLKBUF_X2 inst_16386 ( .A(net_16233), .Z(net_16234) );
AND2_X4 inst_9086 ( .ZN(net_2903), .A2(net_2897), .A1(net_1508) );
CLKBUF_X2 inst_11856 ( .A(net_10667), .Z(net_11704) );
CLKBUF_X2 inst_10233 ( .A(net_10080), .Z(net_10081) );
CLKBUF_X2 inst_10087 ( .A(net_9934), .Z(net_9935) );
INV_X2 inst_6362 ( .ZN(net_2153), .A(net_2152) );
CLKBUF_X2 inst_18377 ( .A(net_18224), .Z(net_18225) );
AOI22_X2 inst_8076 ( .B1(net_8175), .A1(net_7733), .B2(net_6101), .A2(net_6095), .ZN(net_4068) );
CLKBUF_X2 inst_13806 ( .A(net_10369), .Z(net_13654) );
CLKBUF_X2 inst_11009 ( .A(net_10856), .Z(net_10857) );
CLKBUF_X2 inst_10585 ( .A(net_10387), .Z(net_10433) );
XOR2_X2 inst_57 ( .B(net_2969), .A(net_2462), .Z(net_969) );
CLKBUF_X2 inst_15928 ( .A(net_15775), .Z(net_15776) );
CLKBUF_X2 inst_16717 ( .A(net_16564), .Z(net_16565) );
CLKBUF_X2 inst_9312 ( .A(net_9159), .Z(net_9160) );
SDFF_X2 inst_1307 ( .SI(net_7678), .Q(net_7678), .SE(net_2714), .D(net_2702), .CK(net_15296) );
AOI22_X2 inst_7759 ( .B1(net_6987), .A1(net_6947), .A2(net_5443), .B2(net_5442), .ZN(net_5370) );
CLKBUF_X2 inst_10878 ( .A(net_10725), .Z(net_10726) );
AOI22_X2 inst_8565 ( .A1(net_2762), .B2(net_2556), .ZN(net_2298), .A2(net_2030), .B1(net_1750) );
DFF_X1 inst_6789 ( .Q(net_8254), .D(net_4425), .CK(net_18918) );
CLKBUF_X2 inst_16842 ( .A(net_16689), .Z(net_16690) );
CLKBUF_X2 inst_12960 ( .A(net_12807), .Z(net_12808) );
CLKBUF_X2 inst_16925 ( .A(net_16772), .Z(net_16773) );
DFFR_X2 inst_7124 ( .QN(net_7355), .D(net_3065), .CK(net_11622), .RN(x6501) );
AOI222_X1 inst_8616 ( .ZN(net_5032), .A1(net_5031), .A2(net_5030), .B1(net_5029), .B2(net_5028), .C2(net_5027), .C1(net_1518) );
SDFF_X2 inst_851 ( .SI(net_8664), .Q(net_8664), .D(net_3939), .SE(net_3885), .CK(net_12503) );
SDFF_X2 inst_831 ( .SI(net_8630), .Q(net_8630), .D(net_3961), .SE(net_3885), .CK(net_13169) );
CLKBUF_X2 inst_18024 ( .A(net_17871), .Z(net_17872) );
INV_X4 inst_5824 ( .A(net_7506), .ZN(net_4465) );
NAND2_X2 inst_4264 ( .A1(net_7034), .A2(net_5249), .ZN(net_5196) );
CLKBUF_X2 inst_17259 ( .A(net_11439), .Z(net_17107) );
CLKBUF_X2 inst_17668 ( .A(net_9766), .Z(net_17516) );
CLKBUF_X2 inst_11448 ( .A(net_11295), .Z(net_11296) );
NAND2_X2 inst_4430 ( .A1(net_6868), .A2(net_5016), .ZN(net_4997) );
CLKBUF_X2 inst_15007 ( .A(net_11373), .Z(net_14855) );
CLKBUF_X2 inst_11174 ( .A(net_11021), .Z(net_11022) );
SDFF_X2 inst_1497 ( .SI(net_7854), .Q(net_7854), .D(net_2589), .SE(net_2558), .CK(net_18393) );
INV_X4 inst_5706 ( .ZN(net_568), .A(net_263) );
SDFF_X2 inst_1002 ( .D(net_7342), .SI(net_6650), .Q(net_6650), .SE(net_3123), .CK(net_11685) );
CLKBUF_X2 inst_12076 ( .A(net_11923), .Z(net_11924) );
AOI22_X2 inst_8057 ( .B1(net_8139), .A1(net_7901), .A2(net_6098), .ZN(net_6044), .B2(net_4190) );
CLKBUF_X2 inst_13179 ( .A(net_9334), .Z(net_13027) );
SDFF_X2 inst_478 ( .SI(net_8452), .Q(net_8452), .SE(net_3983), .D(net_3981), .CK(net_12461) );
CLKBUF_X2 inst_18985 ( .A(net_18832), .Z(net_18833) );
CLKBUF_X2 inst_18113 ( .A(net_17960), .Z(net_17961) );
AOI222_X1 inst_8630 ( .B2(net_8239), .B1(net_4891), .C2(net_4889), .A1(net_4803), .ZN(net_4767), .C1(net_4465), .A2(net_3384) );
CLKBUF_X2 inst_15832 ( .A(net_15679), .Z(net_15680) );
INV_X4 inst_5666 ( .A(net_6791), .ZN(net_1897) );
CLKBUF_X2 inst_18788 ( .A(net_18635), .Z(net_18636) );
CLKBUF_X2 inst_18219 ( .A(net_18066), .Z(net_18067) );
CLKBUF_X2 inst_13953 ( .A(net_13800), .Z(net_13801) );
CLKBUF_X2 inst_12173 ( .A(net_12020), .Z(net_12021) );
CLKBUF_X2 inst_14126 ( .A(net_13973), .Z(net_13974) );
INV_X4 inst_5378 ( .A(net_1494), .ZN(net_1346) );
INV_X4 inst_5665 ( .A(net_7308), .ZN(net_1258) );
MUX2_X2 inst_4931 ( .A(net_6148), .Z(net_3118), .S(net_2996), .B(net_1051) );
CLKBUF_X2 inst_11540 ( .A(net_11387), .Z(net_11388) );
CLKBUF_X2 inst_15111 ( .A(net_14958), .Z(net_14959) );
DFFR_X2 inst_7334 ( .QN(net_8963), .D(net_2309), .CK(net_14476), .RN(x6501) );
SDFF_X2 inst_799 ( .SI(net_8338), .Q(net_8338), .D(net_3938), .SE(net_3880), .CK(net_10708) );
CLKBUF_X2 inst_12906 ( .A(net_12018), .Z(net_12754) );
NOR2_X2 inst_3481 ( .ZN(net_2243), .A1(net_2242), .A2(net_2241) );
SDFF_X2 inst_738 ( .SI(net_8344), .Q(net_8344), .D(net_3960), .SE(net_3880), .CK(net_13098) );
CLKBUF_X2 inst_13666 ( .A(net_13513), .Z(net_13514) );
INV_X2 inst_6481 ( .A(net_5944), .ZN(x1174) );
CLKBUF_X2 inst_14284 ( .A(net_14131), .Z(net_14132) );
XNOR2_X2 inst_255 ( .B(net_2674), .A(net_2673), .ZN(net_1194) );
SDFFR_X1 inst_2726 ( .SI(net_9038), .Q(net_9038), .D(net_7467), .SE(net_3208), .CK(net_12221), .RN(x6501) );
CLKBUF_X2 inst_10555 ( .A(net_10402), .Z(net_10403) );
SDFFR_X1 inst_2674 ( .SI(net_7539), .SE(net_5043), .CK(net_9714), .RN(x6501), .Q(x4070), .D(x4070) );
CLKBUF_X2 inst_14471 ( .A(net_14002), .Z(net_14319) );
CLKBUF_X2 inst_10390 ( .A(net_10237), .Z(net_10238) );
CLKBUF_X2 inst_10279 ( .A(net_9801), .Z(net_10127) );
HA_X1 inst_6686 ( .A(net_7511), .S(net_3008), .CO(net_3007), .B(net_2974) );
AOI221_X2 inst_8784 ( .C1(net_8979), .B2(net_5538), .C2(net_5456), .ZN(net_5254), .A(net_4930), .B1(net_408) );
SDFF_X2 inst_1113 ( .D(net_7315), .SI(net_6524), .Q(net_6524), .SE(net_3086), .CK(net_9921) );
CLKBUF_X2 inst_12438 ( .A(net_10917), .Z(net_12286) );
NAND2_X2 inst_4206 ( .ZN(net_5289), .A1(net_5050), .A2(net_5049) );
INV_X4 inst_5415 ( .ZN(net_1361), .A(net_863) );
CLKBUF_X2 inst_18398 ( .A(net_18245), .Z(net_18246) );
AOI22_X2 inst_8101 ( .B1(net_8042), .A1(net_8008), .B2(net_6102), .A2(net_6097), .ZN(net_4047) );
SDFFR_X2 inst_2191 ( .SI(net_6485), .Q(net_6485), .SE(net_2933), .D(net_1466), .CK(net_9116), .RN(x6501) );
INV_X4 inst_5296 ( .ZN(net_2318), .A(net_1599) );
SDFF_X2 inst_1127 ( .D(net_7333), .SI(net_6575), .Q(net_6575), .SE(net_3070), .CK(net_9414) );
CLKBUF_X2 inst_12184 ( .A(net_12031), .Z(net_12032) );
SDFF_X2 inst_362 ( .SI(net_8521), .Q(net_8521), .D(net_3980), .SE(net_3979), .CK(net_13378) );
CLKBUF_X2 inst_17013 ( .A(net_13676), .Z(net_16861) );
CLKBUF_X2 inst_19036 ( .A(net_18883), .Z(net_18884) );
XNOR2_X2 inst_306 ( .B(net_7384), .ZN(net_967), .A(net_966) );
AOI222_X1 inst_8662 ( .B1(net_8214), .ZN(net_3601), .A1(net_3600), .A2(net_3599), .B2(net_3598), .C2(net_3597), .C1(net_738) );
CLKBUF_X2 inst_13499 ( .A(net_11635), .Z(net_13347) );
CLKBUF_X2 inst_9460 ( .A(net_9307), .Z(net_9308) );
OAI21_X2 inst_3095 ( .ZN(net_2798), .B2(net_2664), .A(net_2168), .B1(net_1631) );
CLKBUF_X2 inst_9884 ( .A(net_9222), .Z(net_9732) );
SDFF_X2 inst_1715 ( .Q(net_7888), .D(net_7888), .SI(net_2589), .SE(net_2543), .CK(net_15247) );
INV_X2 inst_6396 ( .ZN(net_1165), .A(net_1164) );
CLKBUF_X2 inst_16245 ( .A(net_14787), .Z(net_16093) );
DFFR_X2 inst_7355 ( .Q(net_7329), .CK(net_9534), .D(x13018), .RN(x6501) );
XNOR2_X2 inst_267 ( .B(net_3269), .ZN(net_1096), .A(net_479) );
CLKBUF_X2 inst_16630 ( .A(net_14480), .Z(net_16478) );
CLKBUF_X2 inst_16100 ( .A(net_15947), .Z(net_15948) );
SDFF_X2 inst_716 ( .SI(net_8651), .Q(net_8651), .D(net_3956), .SE(net_3885), .CK(net_10909) );
SDFF_X2 inst_1906 ( .D(net_7270), .SI(net_7007), .Q(net_7007), .SE(net_6277), .CK(net_16802) );
SDFF_X2 inst_792 ( .SI(net_8336), .Q(net_8336), .D(net_3980), .SE(net_3880), .CK(net_10714) );
SDFF_X2 inst_2024 ( .SI(net_7934), .Q(net_7934), .D(net_2710), .SE(net_2461), .CK(net_16452) );
CLKBUF_X2 inst_9984 ( .A(net_9831), .Z(net_9832) );
AND2_X4 inst_9061 ( .A1(net_3320), .A2(net_3305), .ZN(net_3303) );
CLKBUF_X2 inst_16359 ( .A(net_16206), .Z(net_16207) );
CLKBUF_X2 inst_10476 ( .A(net_10261), .Z(net_10324) );
AOI21_X2 inst_8933 ( .B2(net_5843), .ZN(net_5676), .A(net_5675), .B1(x306) );
CLKBUF_X2 inst_16692 ( .A(net_16539), .Z(net_16540) );
SDFFR_X2 inst_2216 ( .Q(net_7473), .D(net_7473), .SE(net_2863), .CK(net_12190), .SI(x13403), .RN(x6501) );
OAI21_X2 inst_2988 ( .B2(net_5912), .ZN(net_5907), .A(net_5801), .B1(net_725) );
CLKBUF_X2 inst_15043 ( .A(net_14890), .Z(net_14891) );
NAND2_X2 inst_4494 ( .A2(net_5538), .ZN(net_4478), .A1(net_428) );
SDFF_X2 inst_1199 ( .D(net_7300), .SI(net_6917), .Q(net_6917), .SE(net_6284), .CK(net_15925) );
CLKBUF_X2 inst_11520 ( .A(net_9400), .Z(net_11368) );
SDFF_X2 inst_1662 ( .SI(net_7755), .Q(net_7755), .D(net_2719), .SE(net_2560), .CK(net_18775) );
DFFR_X1 inst_7508 ( .QN(net_7299), .D(net_1707), .CK(net_18737), .RN(x6501) );
CLKBUF_X2 inst_13240 ( .A(net_13087), .Z(net_13088) );
CLKBUF_X2 inst_11251 ( .A(net_11098), .Z(net_11099) );
SDFF_X2 inst_1285 ( .Q(net_8103), .D(net_8103), .SI(net_2711), .SE(net_2707), .CK(net_14296) );
SDFF_X2 inst_380 ( .SI(net_8399), .Q(net_8399), .SE(net_3969), .D(net_3953), .CK(net_10303) );
CLKBUF_X2 inst_14711 ( .A(net_14558), .Z(net_14559) );
CLKBUF_X2 inst_13508 ( .A(net_13355), .Z(net_13356) );
CLKBUF_X2 inst_18688 ( .A(net_18535), .Z(net_18536) );
DFFR_X1 inst_7423 ( .Q(net_7513), .D(net_4967), .CK(net_13611), .RN(x6501) );
MUX2_X2 inst_4970 ( .B(net_7260), .S(net_2147), .Z(net_1993), .A(net_1492) );
CLKBUF_X2 inst_12583 ( .A(net_12430), .Z(net_12431) );
SDFF_X2 inst_706 ( .SI(net_8628), .Q(net_8628), .SE(net_3984), .D(net_3949), .CK(net_12598) );
CLKBUF_X2 inst_16137 ( .A(net_13640), .Z(net_15985) );
CLKBUF_X2 inst_14692 ( .A(net_14539), .Z(net_14540) );
CLKBUF_X2 inst_10874 ( .A(net_10721), .Z(net_10722) );
CLKBUF_X2 inst_9834 ( .A(net_9681), .Z(net_9682) );
CLKBUF_X2 inst_13366 ( .A(net_13213), .Z(net_13214) );
AOI22_X2 inst_7985 ( .B1(net_8163), .A1(net_7721), .B2(net_6101), .A2(net_6095), .ZN(net_4146) );
NAND2_X2 inst_4734 ( .ZN(net_2584), .A2(net_1586), .A1(net_1118) );
CLKBUF_X2 inst_15033 ( .A(net_14880), .Z(net_14881) );
CLKBUF_X2 inst_13055 ( .A(net_12902), .Z(net_12903) );
XNOR2_X2 inst_110 ( .ZN(net_4705), .A(net_4489), .B(net_940) );
CLKBUF_X2 inst_17927 ( .A(net_17774), .Z(net_17775) );
SDFF_X2 inst_2047 ( .SI(net_7926), .Q(net_7926), .D(net_2590), .SE(net_2461), .CK(net_17648) );
NAND2_X2 inst_4545 ( .ZN(net_3327), .A1(net_3326), .A2(net_3325) );
NAND4_X2 inst_3825 ( .ZN(net_2973), .A1(net_2915), .A2(net_1470), .A3(x2693), .A4(x2633) );
CLKBUF_X2 inst_17740 ( .A(net_17587), .Z(net_17588) );
CLKBUF_X2 inst_16291 ( .A(net_16138), .Z(net_16139) );
AOI22_X2 inst_7876 ( .A1(net_7175), .A2(net_5655), .ZN(net_4565), .B2(net_4564), .B1(net_2499) );
CLKBUF_X2 inst_10842 ( .A(net_10689), .Z(net_10690) );
CLKBUF_X2 inst_11927 ( .A(net_11774), .Z(net_11775) );
AOI22_X2 inst_7846 ( .A2(net_6434), .A1(net_5654), .B2(net_5595), .ZN(net_4662), .B1(net_316) );
CLKBUF_X2 inst_16741 ( .A(net_10321), .Z(net_16589) );
OAI222_X2 inst_2949 ( .A2(net_3889), .B2(net_3888), .C2(net_3887), .ZN(net_3886), .A1(net_2177), .B1(net_1845), .C1(net_508) );
SDFFR_X2 inst_2414 ( .D(net_2690), .SE(net_2313), .SI(net_457), .Q(net_457), .CK(net_13947), .RN(x6501) );
CLKBUF_X2 inst_18224 ( .A(net_17024), .Z(net_18072) );
CLKBUF_X2 inst_10429 ( .A(net_10276), .Z(net_10277) );
CLKBUF_X2 inst_11132 ( .A(net_10979), .Z(net_10980) );
AOI22_X2 inst_7901 ( .A2(net_5538), .ZN(net_4527), .B1(net_4526), .B2(net_4388), .A1(net_411) );
CLKBUF_X2 inst_15189 ( .A(net_14287), .Z(net_15037) );
DFFR_X2 inst_6981 ( .QN(net_5964), .D(net_5903), .CK(net_9282), .RN(x6501) );
CLKBUF_X2 inst_11695 ( .A(net_10714), .Z(net_11543) );
CLKBUF_X2 inst_14648 ( .A(net_14495), .Z(net_14496) );
DFFR_X2 inst_7316 ( .D(net_8285), .QN(net_8281), .CK(net_12225), .RN(x6501) );
CLKBUF_X2 inst_16619 ( .A(net_16466), .Z(net_16467) );
CLKBUF_X2 inst_14440 ( .A(net_14287), .Z(net_14288) );
SDFF_X2 inst_889 ( .Q(net_8558), .D(net_8558), .SI(net_3980), .SE(net_3878), .CK(net_13303) );
AOI21_X2 inst_8935 ( .B2(net_5871), .ZN(net_5669), .A(net_5668), .B1(net_2744) );
AOI22_X2 inst_8533 ( .B1(net_6724), .A1(net_6691), .B2(net_6202), .A2(net_3520), .ZN(net_3407) );
CLKBUF_X2 inst_16302 ( .A(net_16149), .Z(net_16150) );
CLKBUF_X2 inst_12457 ( .A(net_12304), .Z(net_12305) );
INV_X4 inst_5188 ( .ZN(net_2915), .A(net_2747) );
SDFFR_X2 inst_2379 ( .SE(net_2260), .Q(net_317), .D(net_317), .CK(net_9295), .RN(x6501), .SI(x3258) );
CLKBUF_X2 inst_10358 ( .A(net_10205), .Z(net_10206) );
AOI221_X2 inst_8774 ( .B1(net_5268), .C2(net_5267), .ZN(net_5265), .A(net_4915), .B2(net_4626), .C1(net_172) );
CLKBUF_X2 inst_11754 ( .A(net_11359), .Z(net_11602) );
CLKBUF_X2 inst_11244 ( .A(net_10943), .Z(net_11092) );
CLKBUF_X2 inst_15047 ( .A(net_14894), .Z(net_14895) );
CLKBUF_X2 inst_16275 ( .A(net_16122), .Z(net_16123) );
CLKBUF_X2 inst_10382 ( .A(net_10229), .Z(net_10230) );
MUX2_X2 inst_4916 ( .B(net_6320), .Z(net_5526), .A(net_5525), .S(net_5522) );
AOI22_X2 inst_8149 ( .B1(net_8086), .A1(net_7746), .B2(net_6108), .A2(net_6096), .ZN(net_4003) );
NOR2_X2 inst_3571 ( .A1(net_6753), .A2(net_6752), .ZN(net_2901) );
CLKBUF_X2 inst_15757 ( .A(net_15604), .Z(net_15605) );
INV_X4 inst_6132 ( .A(net_6410), .ZN(net_1316) );
SDFF_X2 inst_1190 ( .D(net_7328), .SI(net_6570), .Q(net_6570), .SE(net_3070), .CK(net_11746) );
SDFF_X2 inst_444 ( .Q(net_8773), .D(net_8773), .SE(net_3982), .SI(net_3950), .CK(net_10584) );
AOI221_X2 inst_8865 ( .ZN(net_2986), .C2(net_2133), .C1(net_2008), .B1(net_1910), .A(net_1669), .B2(net_1475) );
DFFR_X1 inst_7489 ( .QN(net_7632), .D(net_3903), .CK(net_11266), .RN(x6501) );
AOI22_X2 inst_8246 ( .B1(net_8798), .A1(net_8539), .A2(net_3861), .B2(net_3860), .ZN(net_3791) );
CLKBUF_X2 inst_12816 ( .A(net_12663), .Z(net_12664) );
AND2_X4 inst_9064 ( .ZN(net_6110), .A2(net_3249), .A1(net_3248) );
CLKBUF_X2 inst_10033 ( .A(net_9880), .Z(net_9881) );
CLKBUF_X2 inst_14196 ( .A(net_12485), .Z(net_14044) );
AOI221_X4 inst_8705 ( .C1(net_8193), .B1(net_7683), .C2(net_6099), .ZN(net_6033), .B2(net_4399), .A(net_4306) );
CLKBUF_X2 inst_11720 ( .A(net_11567), .Z(net_11568) );
CLKBUF_X2 inst_18612 ( .A(net_11570), .Z(net_18460) );
INV_X4 inst_5833 ( .A(net_6355), .ZN(net_727) );
CLKBUF_X2 inst_12047 ( .A(net_11894), .Z(net_11895) );
XNOR2_X2 inst_119 ( .A(net_3022), .ZN(net_3001), .B(net_3000) );
OAI211_X2 inst_3181 ( .B(net_6124), .ZN(net_5598), .C2(net_5533), .A(net_2946), .C1(net_2842) );
SDFF_X2 inst_939 ( .SI(net_7318), .Q(net_6659), .D(net_6659), .SE(net_3126), .CK(net_12150) );
CLKBUF_X2 inst_9722 ( .A(net_9569), .Z(net_9570) );
CLKBUF_X2 inst_17912 ( .A(net_15576), .Z(net_17760) );
CLKBUF_X2 inst_10770 ( .A(net_9081), .Z(net_10618) );
CLKBUF_X2 inst_18609 ( .A(net_18456), .Z(net_18457) );
AOI22_X2 inst_8205 ( .B1(net_8793), .A1(net_8534), .A2(net_3861), .B2(net_3860), .ZN(net_3831) );
CLKBUF_X2 inst_15389 ( .A(net_15236), .Z(net_15237) );
SDFF_X2 inst_1019 ( .SI(net_7334), .Q(net_6675), .D(net_6675), .SE(net_3126), .CK(net_12022) );
CLKBUF_X2 inst_17364 ( .A(net_17211), .Z(net_17212) );
CLKBUF_X2 inst_13490 ( .A(net_13337), .Z(net_13338) );
CLKBUF_X2 inst_16748 ( .A(net_16595), .Z(net_16596) );
CLKBUF_X2 inst_15672 ( .A(net_15519), .Z(net_15520) );
SDFF_X2 inst_1827 ( .D(net_7281), .SI(net_6858), .Q(net_6858), .SE(net_6282), .CK(net_19004) );
CLKBUF_X2 inst_10830 ( .A(net_9851), .Z(net_10678) );
SDFF_X2 inst_742 ( .Q(net_8805), .D(net_8805), .SI(net_3941), .SE(net_3879), .CK(net_12874) );
CLKBUF_X2 inst_13372 ( .A(net_9522), .Z(net_13220) );
NAND2_X2 inst_4481 ( .A2(net_5267), .ZN(net_4497), .A1(net_181) );
CLKBUF_X2 inst_17888 ( .A(net_17735), .Z(net_17736) );
CLKBUF_X2 inst_13545 ( .A(net_12937), .Z(net_13393) );
DFFR_X2 inst_7345 ( .Q(net_7332), .CK(net_11661), .D(x12991), .RN(x6501) );
INV_X4 inst_5289 ( .ZN(net_1782), .A(net_1379) );
AND2_X4 inst_9121 ( .A2(net_7209), .ZN(net_2085), .A1(net_1083) );
SDFF_X2 inst_1955 ( .D(net_7297), .SI(net_6914), .Q(net_6914), .SE(net_6284), .CK(net_18178) );
CLKBUF_X2 inst_18287 ( .A(net_18134), .Z(net_18135) );
NOR2_X2 inst_3618 ( .A2(net_7526), .A1(net_7524), .ZN(net_1617) );
CLKBUF_X2 inst_17533 ( .A(net_17380), .Z(net_17381) );
CLKBUF_X2 inst_14807 ( .A(net_14654), .Z(net_14655) );
CLKBUF_X2 inst_14430 ( .A(net_14277), .Z(net_14278) );
CLKBUF_X2 inst_14945 ( .A(net_11750), .Z(net_14793) );
AND2_X2 inst_9181 ( .A2(net_6093), .ZN(net_2781), .A1(net_2028) );
CLKBUF_X2 inst_9781 ( .A(net_9483), .Z(net_9629) );
SDFFR_X1 inst_2704 ( .SI(net_7536), .SE(net_5043), .CK(net_9683), .RN(x6501), .Q(x4104), .D(x4104) );
AOI22_X2 inst_8349 ( .B1(net_8812), .A1(net_8553), .A2(net_3861), .B2(net_3860), .ZN(net_3699) );
CLKBUF_X2 inst_11461 ( .A(net_11308), .Z(net_11309) );
CLKBUF_X2 inst_18828 ( .A(net_18675), .Z(net_18676) );
INV_X4 inst_5924 ( .A(net_6290), .ZN(net_2727) );
CLKBUF_X2 inst_14551 ( .A(net_9930), .Z(net_14399) );
CLKBUF_X2 inst_13327 ( .A(net_13174), .Z(net_13175) );
CLKBUF_X2 inst_9508 ( .A(net_9355), .Z(net_9356) );
CLKBUF_X2 inst_16355 ( .A(net_16202), .Z(net_16203) );
CLKBUF_X2 inst_9701 ( .A(net_9215), .Z(net_9549) );
INV_X4 inst_5473 ( .A(net_1622), .ZN(net_746) );
CLKBUF_X2 inst_15014 ( .A(net_14861), .Z(net_14862) );
CLKBUF_X2 inst_18290 ( .A(net_18137), .Z(net_18138) );
NAND2_X2 inst_4817 ( .ZN(net_1247), .A1(net_803), .A2(net_730) );
NAND2_X2 inst_4456 ( .ZN(net_4949), .A2(net_4833), .A1(net_4500) );
MUX2_X2 inst_4926 ( .Z(net_3553), .S(net_3552), .B(net_999), .A(net_976) );
DFF_X1 inst_6846 ( .QN(net_6425), .D(net_3635), .CK(net_17959) );
CLKBUF_X2 inst_13840 ( .A(net_13687), .Z(net_13688) );
NAND2_X2 inst_4571 ( .A1(net_8255), .ZN(net_6084), .A2(net_3028) );
INV_X4 inst_5111 ( .ZN(net_4945), .A(net_4878) );
NAND3_X2 inst_3928 ( .ZN(net_5591), .A3(net_5465), .A2(net_4491), .A1(net_4490) );
CLKBUF_X2 inst_12212 ( .A(net_12059), .Z(net_12060) );
CLKBUF_X2 inst_11849 ( .A(net_10251), .Z(net_11697) );
NAND2_X4 inst_4017 ( .A2(net_6796), .A1(net_6271), .ZN(net_4375) );
DFFR_X2 inst_7121 ( .QN(net_7601), .D(net_3078), .CK(net_9793), .RN(x6501) );
CLKBUF_X2 inst_19054 ( .A(net_18901), .Z(net_18902) );
CLKBUF_X2 inst_16917 ( .A(net_16764), .Z(net_16765) );
CLKBUF_X2 inst_18723 ( .A(net_18570), .Z(net_18571) );
INV_X4 inst_5135 ( .ZN(net_4221), .A(net_3552) );
CLKBUF_X2 inst_17216 ( .A(net_11501), .Z(net_17064) );
CLKBUF_X2 inst_12879 ( .A(net_12726), .Z(net_12727) );
CLKBUF_X2 inst_13050 ( .A(net_12527), .Z(net_12898) );
INV_X4 inst_5760 ( .A(net_7578), .ZN(net_559) );
DFFR_X1 inst_7556 ( .D(net_7303), .QN(net_6416), .CK(net_9664), .RN(x6501) );
CLKBUF_X2 inst_11513 ( .A(net_10100), .Z(net_11361) );
DFFR_X2 inst_7037 ( .QN(net_7503), .D(net_4974), .CK(net_14506), .RN(x6501) );
DFFR_X2 inst_7294 ( .Q(net_6411), .D(net_1079), .CK(net_17990), .RN(x6501) );
INV_X4 inst_5095 ( .ZN(net_5702), .A(net_5676) );
CLKBUF_X2 inst_14591 ( .A(net_14438), .Z(net_14439) );
CLKBUF_X2 inst_17760 ( .A(net_17607), .Z(net_17608) );
CLKBUF_X2 inst_17905 ( .A(net_17752), .Z(net_17753) );
CLKBUF_X2 inst_18636 ( .A(net_18483), .Z(net_18484) );
SDFF_X2 inst_426 ( .Q(net_8753), .D(net_8753), .SE(net_3982), .SI(net_3945), .CK(net_13065) );
INV_X4 inst_6035 ( .A(net_7350), .ZN(net_3079) );
CLKBUF_X2 inst_13856 ( .A(net_13703), .Z(net_13704) );
NAND2_X2 inst_4302 ( .A1(net_7133), .A2(net_5166), .ZN(net_5155) );
CLKBUF_X2 inst_11654 ( .A(net_11501), .Z(net_11502) );
CLKBUF_X2 inst_11068 ( .A(net_10915), .Z(net_10916) );
AOI22_X2 inst_8092 ( .B1(net_8143), .A1(net_7905), .A2(net_6098), .ZN(net_6052), .B2(net_4190) );
INV_X2 inst_6560 ( .A(net_7566), .ZN(net_3132) );
INV_X2 inst_6341 ( .ZN(net_2591), .A(net_2527) );
CLKBUF_X2 inst_16875 ( .A(net_16722), .Z(net_16723) );
CLKBUF_X2 inst_11163 ( .A(net_11010), .Z(net_11011) );
AOI22_X2 inst_8544 ( .B1(net_6528), .A1(net_6495), .A2(net_6137), .B2(net_6104), .ZN(net_3396) );
CLKBUF_X2 inst_9247 ( .A(net_9094), .Z(net_9095) );
CLKBUF_X2 inst_9904 ( .A(net_9751), .Z(net_9752) );
CLKBUF_X2 inst_15182 ( .A(net_15029), .Z(net_15030) );
CLKBUF_X2 inst_12558 ( .A(net_12405), .Z(net_12406) );
AOI22_X2 inst_8136 ( .B1(net_8118), .A1(net_7880), .A2(net_6098), .B2(net_4190), .ZN(net_4014) );
CLKBUF_X2 inst_15645 ( .A(net_15492), .Z(net_15493) );
CLKBUF_X2 inst_19055 ( .A(net_9512), .Z(net_18903) );
NAND2_X2 inst_4211 ( .A1(net_6880), .ZN(net_5251), .A2(net_5247) );
SDFF_X2 inst_1745 ( .Q(net_7901), .D(net_7901), .SI(net_2639), .SE(net_2543), .CK(net_17116) );
NAND4_X2 inst_3831 ( .A1(net_9052), .A4(net_6250), .A3(net_2946), .A2(net_2532), .ZN(net_2348) );
SDFFS_X2 inst_2079 ( .SI(net_7384), .SE(net_2795), .Q(net_173), .D(net_173), .CK(net_17493), .SN(x6501) );
CLKBUF_X2 inst_10534 ( .A(net_10381), .Z(net_10382) );
CLKBUF_X2 inst_15506 ( .A(net_15353), .Z(net_15354) );
DFF_X1 inst_6819 ( .QN(net_8232), .D(net_4449), .CK(net_17208) );
CLKBUF_X2 inst_19106 ( .A(net_16106), .Z(net_18954) );
CLKBUF_X2 inst_18057 ( .A(net_17904), .Z(net_17905) );
CLKBUF_X2 inst_14883 ( .A(net_14730), .Z(net_14731) );
CLKBUF_X2 inst_9299 ( .A(net_9146), .Z(net_9147) );
CLKBUF_X2 inst_19120 ( .A(net_18967), .Z(net_18968) );
CLKBUF_X2 inst_14053 ( .A(net_12929), .Z(net_13901) );
INV_X2 inst_6554 ( .A(net_8952), .ZN(net_789) );
INV_X4 inst_5615 ( .A(net_8919), .ZN(net_4526) );
CLKBUF_X2 inst_14729 ( .A(net_14576), .Z(net_14577) );
CLKBUF_X2 inst_12081 ( .A(net_10374), .Z(net_11929) );
SDFFR_X2 inst_2596 ( .Q(net_7303), .D(net_7303), .SE(net_1578), .SI(net_1576), .CK(net_15144), .RN(x6501) );
CLKBUF_X2 inst_18575 ( .A(net_18422), .Z(net_18423) );
INV_X2 inst_6599 ( .A(net_6147), .ZN(net_6146) );
INV_X2 inst_6242 ( .ZN(net_4894), .A(net_4797) );
AOI22_X2 inst_8579 ( .B1(net_2569), .A2(net_1588), .B2(net_1517), .ZN(net_1516), .A1(net_1515) );
OAI21_X2 inst_3022 ( .ZN(net_4976), .A(net_4826), .B2(net_4382), .B1(net_262) );
CLKBUF_X2 inst_12133 ( .A(net_11980), .Z(net_11981) );
SDFF_X2 inst_680 ( .Q(net_8697), .D(net_8697), .SI(net_3940), .SE(net_3935), .CK(net_10349) );
INV_X2 inst_6575 ( .ZN(net_802), .A(net_227) );
CLKBUF_X2 inst_10323 ( .A(net_9249), .Z(net_10171) );
NOR3_X2 inst_3299 ( .ZN(net_1852), .A2(net_1571), .A3(net_1566), .A1(net_1305) );
CLKBUF_X2 inst_16565 ( .A(net_10173), .Z(net_16413) );
AOI22_X2 inst_7820 ( .A2(net_8253), .B1(net_5029), .ZN(net_4730), .A1(net_4729), .B2(net_4728) );
DFFR_X2 inst_7065 ( .QN(net_7486), .D(net_4268), .CK(net_11251), .RN(x6501) );
CLKBUF_X2 inst_15717 ( .A(net_13220), .Z(net_15565) );
DFFR_X1 inst_7551 ( .QN(net_5950), .D(net_918), .CK(net_11631), .RN(x6501) );
CLKBUF_X2 inst_12697 ( .A(net_12544), .Z(net_12545) );
NOR2_X2 inst_3567 ( .A2(net_6142), .A1(net_6139), .ZN(net_1180) );
CLKBUF_X2 inst_16223 ( .A(net_16070), .Z(net_16071) );
SDFF_X2 inst_414 ( .SI(net_8328), .Q(net_8328), .SE(net_3978), .D(net_3951), .CK(net_10610) );
CLKBUF_X2 inst_18261 ( .A(net_17797), .Z(net_18109) );
SDFF_X2 inst_531 ( .Q(net_8888), .D(net_8888), .SI(net_3948), .SE(net_3936), .CK(net_13480) );
CLKBUF_X2 inst_9315 ( .A(net_9162), .Z(net_9163) );
SDFF_X2 inst_1952 ( .D(net_7263), .SI(net_6920), .Q(net_6920), .SE(net_6281), .CK(net_14319) );
AOI221_X2 inst_8827 ( .C1(net_8161), .B1(net_7719), .C2(net_6101), .B2(net_6095), .ZN(net_6003), .A(net_4304) );
INV_X4 inst_6060 ( .A(net_6350), .ZN(net_493) );
INV_X8 inst_5023 ( .ZN(net_4365), .A(net_3355) );
INV_X4 inst_5617 ( .A(net_8920), .ZN(net_2616) );
NAND4_X2 inst_3698 ( .ZN(net_4439), .A4(net_4340), .A1(net_3775), .A2(net_3774), .A3(net_3773) );
NAND2_X2 inst_4155 ( .ZN(net_5360), .A1(net_5101), .A2(net_5100) );
DFFS_X1 inst_6962 ( .D(net_1143), .CK(net_16326), .SN(x6501), .Q(x919) );
INV_X4 inst_5118 ( .A(net_8225), .ZN(net_4847) );
CLKBUF_X2 inst_14223 ( .A(net_14070), .Z(net_14071) );
CLKBUF_X2 inst_9686 ( .A(net_9533), .Z(net_9534) );
CLKBUF_X2 inst_15102 ( .A(net_14949), .Z(net_14950) );
CLKBUF_X2 inst_10208 ( .A(net_10055), .Z(net_10056) );
CLKBUF_X2 inst_16944 ( .A(net_16791), .Z(net_16792) );
CLKBUF_X2 inst_17771 ( .A(net_17618), .Z(net_17619) );
CLKBUF_X2 inst_10699 ( .A(net_10546), .Z(net_10547) );
INV_X4 inst_5338 ( .ZN(net_1452), .A(net_1317) );
SDFF_X2 inst_570 ( .Q(net_8816), .D(net_8816), .SE(net_3964), .SI(net_3943), .CK(net_10737) );
SDFF_X2 inst_1570 ( .SI(net_7713), .Q(net_7713), .D(net_2573), .SE(net_2559), .CK(net_18048) );
CLKBUF_X2 inst_14697 ( .A(net_14544), .Z(net_14545) );
CLKBUF_X2 inst_16424 ( .A(net_16271), .Z(net_16272) );
CLKBUF_X2 inst_12055 ( .A(net_11902), .Z(net_11903) );
SDFF_X2 inst_1612 ( .Q(net_8119), .D(net_8119), .SI(net_2658), .SE(net_2541), .CK(net_15516) );
NAND2_X2 inst_4645 ( .ZN(net_2347), .A1(net_2346), .A2(net_2339) );
CLKBUF_X2 inst_16054 ( .A(net_13780), .Z(net_15902) );
CLKBUF_X2 inst_12545 ( .A(net_12392), .Z(net_12393) );
CLKBUF_X2 inst_15649 ( .A(net_14698), .Z(net_15497) );
CLKBUF_X2 inst_17295 ( .A(net_17142), .Z(net_17143) );
CLKBUF_X2 inst_11419 ( .A(net_10209), .Z(net_11267) );
NAND4_X2 inst_3718 ( .ZN(net_4419), .A4(net_4328), .A1(net_3649), .A2(net_3648), .A3(net_3647) );
CLKBUF_X2 inst_12592 ( .A(net_12439), .Z(net_12440) );
OAI21_X2 inst_3077 ( .ZN(net_3881), .B2(net_3552), .B1(net_3278), .A(net_873) );
CLKBUF_X2 inst_18675 ( .A(net_9696), .Z(net_18523) );
CLKBUF_X2 inst_15905 ( .A(net_15752), .Z(net_15753) );
CLKBUF_X2 inst_12599 ( .A(net_12446), .Z(net_12447) );
INV_X4 inst_5224 ( .A(net_2453), .ZN(net_2280) );
AOI22_X2 inst_8099 ( .B1(net_8144), .A1(net_7906), .A2(net_6098), .ZN(net_6059), .B2(net_4190) );
CLKBUF_X2 inst_9566 ( .A(net_9413), .Z(net_9414) );
SDFF_X2 inst_1423 ( .SI(net_7279), .Q(net_7056), .D(net_7056), .SE(net_6280), .CK(net_19044) );
SDFF_X2 inst_1034 ( .SI(net_7327), .Q(net_6734), .D(net_6734), .SE(net_3124), .CK(net_9095) );
CLKBUF_X2 inst_15448 ( .A(net_15295), .Z(net_15296) );
CLKBUF_X2 inst_9855 ( .A(net_9702), .Z(net_9703) );
SDFF_X2 inst_1207 ( .Q(net_8101), .D(net_8101), .SI(net_2749), .SE(net_2707), .CK(net_13807) );
CLKBUF_X2 inst_14492 ( .A(net_9328), .Z(net_14340) );
SDFF_X2 inst_613 ( .SI(net_8375), .Q(net_8375), .SE(net_3969), .D(net_3938), .CK(net_13048) );
CLKBUF_X2 inst_9945 ( .A(net_9792), .Z(net_9793) );
NAND2_X2 inst_4275 ( .A1(net_6919), .A2(net_5247), .ZN(net_5185) );
AOI222_X1 inst_8694 ( .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3206), .C1(net_3205), .B1(net_3141), .A2(net_3017) );
INV_X2 inst_6444 ( .ZN(net_869), .A(net_607) );
SDFF_X2 inst_483 ( .SI(net_8605), .Q(net_8605), .SE(net_3984), .D(net_3945), .CK(net_13141) );
CLKBUF_X2 inst_16186 ( .A(net_11284), .Z(net_16034) );
MUX2_X2 inst_5005 ( .A(net_9018), .B(net_6203), .Z(net_3977), .S(net_622) );
CLKBUF_X2 inst_9907 ( .A(net_9754), .Z(net_9755) );
XNOR2_X2 inst_259 ( .ZN(net_1187), .A(net_1186), .B(net_846) );
CLKBUF_X2 inst_17652 ( .A(net_17499), .Z(net_17500) );
DFF_X1 inst_6845 ( .QN(net_6424), .D(net_3610), .CK(net_17962) );
CLKBUF_X2 inst_17659 ( .A(net_17506), .Z(net_17507) );
DFF_X1 inst_6812 ( .Q(net_8253), .D(net_4426), .CK(net_17588) );
NAND2_X2 inst_4707 ( .A1(net_7368), .A2(net_1885), .ZN(net_1859) );
NAND2_X2 inst_4846 ( .ZN(net_906), .A1(net_677), .A2(net_524) );
AOI222_X1 inst_8621 ( .A2(net_8225), .A1(net_4891), .B2(net_4889), .C2(net_4888), .ZN(net_4885), .B1(net_4884), .C1(net_3110) );
CLKBUF_X2 inst_13197 ( .A(net_13044), .Z(net_13045) );
CLKBUF_X2 inst_10517 ( .A(net_10364), .Z(net_10365) );
CLKBUF_X2 inst_10686 ( .A(net_10533), .Z(net_10534) );
CLKBUF_X2 inst_16217 ( .A(net_10637), .Z(net_16065) );
SDFF_X2 inst_894 ( .Q(net_8571), .D(net_8571), .SI(net_3973), .SE(net_3878), .CK(net_12327) );
CLKBUF_X2 inst_19083 ( .A(net_18930), .Z(net_18931) );
SDFFR_X2 inst_2425 ( .D(net_2676), .SE(net_2313), .SI(net_475), .Q(net_475), .CK(net_16902), .RN(x6501) );
CLKBUF_X2 inst_16645 ( .A(net_16492), .Z(net_16493) );
SDFF_X2 inst_994 ( .D(net_7332), .SI(net_6640), .Q(net_6640), .SE(net_3123), .CK(net_9077) );
CLKBUF_X2 inst_9803 ( .A(net_9644), .Z(net_9651) );
SDFF_X2 inst_1879 ( .D(net_7287), .SI(net_6984), .Q(net_6984), .SE(net_6283), .CK(net_14877) );
SDFF_X2 inst_1863 ( .D(net_7296), .SI(net_6873), .Q(net_6873), .SE(net_6282), .CK(net_15412) );
SDFFR_X2 inst_2135 ( .SI(net_7203), .Q(net_7203), .D(net_6454), .SE(net_4362), .CK(net_13728), .RN(x6501) );
CLKBUF_X2 inst_17439 ( .A(net_17286), .Z(net_17287) );
CLKBUF_X2 inst_14082 ( .A(net_13929), .Z(net_13930) );
SDFF_X2 inst_764 ( .Q(net_8807), .D(net_8807), .SI(net_3952), .SE(net_3879), .CK(net_12869) );
CLKBUF_X2 inst_17764 ( .A(net_17611), .Z(net_17612) );
CLKBUF_X2 inst_10961 ( .A(net_10020), .Z(net_10809) );
CLKBUF_X2 inst_12015 ( .A(net_11862), .Z(net_11863) );
SDFF_X2 inst_1547 ( .Q(net_8003), .D(net_8003), .SI(net_2639), .SE(net_2542), .CK(net_16497) );
CLKBUF_X2 inst_11745 ( .A(net_11592), .Z(net_11593) );
SDFFR_X2 inst_2369 ( .D(net_7366), .SI(net_2701), .SE(net_2345), .QN(net_267), .CK(net_16118), .RN(x6501) );
CLKBUF_X2 inst_18482 ( .A(net_16019), .Z(net_18330) );
INV_X4 inst_6105 ( .A(net_7377), .ZN(net_1117) );
SDFF_X2 inst_1274 ( .Q(net_7839), .D(net_7839), .SE(net_2730), .SI(net_2703), .CK(net_14029) );
NAND4_X2 inst_3838 ( .ZN(net_2287), .A2(net_2047), .A4(net_2046), .A3(net_1863), .A1(net_1689) );
CLKBUF_X2 inst_16444 ( .A(net_16291), .Z(net_16292) );
INV_X4 inst_5495 ( .ZN(net_717), .A(net_716) );
INV_X4 inst_5326 ( .A(net_1380), .ZN(net_1355) );
CLKBUF_X2 inst_14847 ( .A(net_14694), .Z(net_14695) );
DFFR_X2 inst_7237 ( .QN(net_6834), .D(net_2195), .CK(net_18723), .RN(x6501) );
OR2_X4 inst_2831 ( .ZN(net_3031), .A2(net_2999), .A1(net_522) );
CLKBUF_X2 inst_12785 ( .A(net_12632), .Z(net_12633) );
SDFF_X2 inst_1300 ( .Q(net_8094), .D(net_8094), .SE(net_2707), .SI(net_2575), .CK(net_16008) );
CLKBUF_X2 inst_12022 ( .A(net_11869), .Z(net_11870) );
INV_X4 inst_5317 ( .ZN(net_1814), .A(net_1813) );
CLKBUF_X2 inst_13698 ( .A(net_13545), .Z(net_13546) );
CLKBUF_X2 inst_13693 ( .A(net_13540), .Z(net_13541) );
DFFR_X2 inst_7309 ( .D(net_290), .QN(net_149), .CK(net_9640), .RN(x6501) );
CLKBUF_X2 inst_15284 ( .A(net_13370), .Z(net_15132) );
SDFFR_X2 inst_2279 ( .SI(net_7392), .SE(net_2789), .Q(net_251), .D(net_251), .CK(net_17764), .RN(x6501) );
CLKBUF_X2 inst_12572 ( .A(net_9128), .Z(net_12420) );
SDFF_X2 inst_2038 ( .SI(net_7783), .Q(net_7783), .D(net_2706), .SE(net_2459), .CK(net_18834) );
SDFF_X2 inst_2044 ( .SI(net_7931), .Q(net_7931), .D(net_2749), .SE(net_2461), .CK(net_16446) );
CLKBUF_X2 inst_19109 ( .A(net_18956), .Z(net_18957) );
AOI22_X2 inst_7833 ( .A2(net_5535), .B2(net_5260), .ZN(net_4688), .B1(net_3111), .A1(net_460) );
CLKBUF_X2 inst_15820 ( .A(net_15667), .Z(net_15668) );
CLKBUF_X2 inst_15289 ( .A(net_12340), .Z(net_15137) );
CLKBUF_X2 inst_13630 ( .A(net_11480), .Z(net_13478) );
INV_X2 inst_6249 ( .ZN(net_4857), .A(net_4745) );
CLKBUF_X2 inst_15245 ( .A(net_12445), .Z(net_15093) );
CLKBUF_X2 inst_13711 ( .A(net_13558), .Z(net_13559) );
INV_X2 inst_6610 ( .A(net_6200), .ZN(net_6198) );
SDFFR_X2 inst_2493 ( .Q(net_8994), .D(net_8994), .SI(net_2604), .SE(net_2562), .CK(net_14801), .RN(x6501) );
SDFF_X2 inst_511 ( .Q(net_8864), .D(net_8864), .SI(net_3945), .SE(net_3936), .CK(net_11096) );
CLKBUF_X2 inst_9593 ( .A(net_9239), .Z(net_9441) );
AOI222_X1 inst_8665 ( .A1(net_7653), .C1(net_7649), .A2(net_3599), .B2(net_3598), .C2(net_3597), .ZN(net_3593), .B1(net_1471) );
CLKBUF_X2 inst_14720 ( .A(net_14567), .Z(net_14568) );
SDFFR_X1 inst_2645 ( .D(net_6768), .SE(net_4506), .CK(net_9251), .RN(x6501), .SI(x1829), .Q(x1829) );
SDFF_X2 inst_1164 ( .SI(net_7318), .Q(net_6593), .D(net_6593), .SE(net_3069), .CK(net_9900) );
CLKBUF_X2 inst_18369 ( .A(net_10686), .Z(net_18217) );
OAI21_X2 inst_3112 ( .ZN(net_2436), .A(net_2435), .B2(net_2385), .B1(net_1859) );
CLKBUF_X2 inst_14025 ( .A(net_13872), .Z(net_13873) );
CLKBUF_X2 inst_11410 ( .A(net_11257), .Z(net_11258) );
CLKBUF_X2 inst_15994 ( .A(net_12489), .Z(net_15842) );
DFFR_X2 inst_7276 ( .QN(net_6341), .D(net_6339), .CK(net_16929), .RN(x6501) );
CLKBUF_X2 inst_15340 ( .A(net_13400), .Z(net_15188) );
CLKBUF_X2 inst_15501 ( .A(net_15348), .Z(net_15349) );
CLKBUF_X2 inst_14613 ( .A(net_11847), .Z(net_14461) );
CLKBUF_X2 inst_18742 ( .A(net_18589), .Z(net_18590) );
CLKBUF_X2 inst_11416 ( .A(net_11263), .Z(net_11264) );
CLKBUF_X2 inst_14596 ( .A(net_10330), .Z(net_14444) );
SDFF_X2 inst_1242 ( .Q(net_7975), .D(net_7975), .SE(net_2755), .SI(net_2703), .CK(net_16879) );
CLKBUF_X2 inst_16558 ( .A(net_16405), .Z(net_16406) );
CLKBUF_X2 inst_14915 ( .A(net_14762), .Z(net_14763) );
CLKBUF_X2 inst_14578 ( .A(net_14425), .Z(net_14426) );
CLKBUF_X2 inst_18849 ( .A(net_18696), .Z(net_18697) );
CLKBUF_X2 inst_17838 ( .A(net_15683), .Z(net_17686) );
CLKBUF_X2 inst_13363 ( .A(net_11866), .Z(net_13211) );
AOI22_X2 inst_8362 ( .B1(net_8777), .A1(net_8407), .A2(net_3867), .B2(net_3866), .ZN(net_3686) );
SDFF_X2 inst_388 ( .Q(net_8848), .D(net_8848), .SI(net_3976), .SE(net_3964), .CK(net_12561) );
CLKBUF_X2 inst_12374 ( .A(net_9714), .Z(net_12222) );
CLKBUF_X2 inst_15119 ( .A(net_14966), .Z(net_14967) );
SDFF_X2 inst_489 ( .SI(net_8594), .Q(net_8594), .SE(net_3984), .D(net_3943), .CK(net_13139) );
CLKBUF_X2 inst_9278 ( .A(net_9061), .Z(net_9126) );
INV_X4 inst_5502 ( .A(net_1236), .ZN(net_801) );
DFFR_X2 inst_7153 ( .QN(net_7219), .D(net_2862), .CK(net_16159), .RN(x6501) );
NOR2_X1 inst_3622 ( .A2(net_6325), .ZN(net_1505), .A1(net_826) );
CLKBUF_X2 inst_18041 ( .A(net_13117), .Z(net_17889) );
CLKBUF_X2 inst_11625 ( .A(net_11472), .Z(net_11473) );
XOR2_X2 inst_39 ( .B(net_3127), .Z(net_1094), .A(net_1093) );
SDFFR_X2 inst_2627 ( .Q(net_7378), .D(net_7378), .SE(net_1136), .CK(net_9059), .RN(x6501), .SI(x4757) );
AOI21_X2 inst_8987 ( .ZN(net_1891), .A(net_1821), .B2(net_1819), .B1(net_1653) );
OAI21_X2 inst_3173 ( .ZN(net_5981), .A(net_3003), .B1(net_2848), .B2(net_1797) );
XNOR2_X2 inst_125 ( .ZN(net_2878), .B(net_2829), .A(net_2828) );
NAND2_X2 inst_4770 ( .ZN(net_1923), .A2(net_1662), .A1(net_484) );
CLKBUF_X2 inst_15517 ( .A(net_15364), .Z(net_15365) );
CLKBUF_X2 inst_17134 ( .A(net_16981), .Z(net_16982) );
CLKBUF_X2 inst_15233 ( .A(net_15080), .Z(net_15081) );
CLKBUF_X2 inst_11919 ( .A(net_11766), .Z(net_11767) );
CLKBUF_X2 inst_14753 ( .A(net_14600), .Z(net_14601) );
CLKBUF_X2 inst_17557 ( .A(net_17404), .Z(net_17405) );
SDFF_X2 inst_430 ( .Q(net_8758), .D(net_8758), .SE(net_3982), .SI(net_3967), .CK(net_13063) );
CLKBUF_X2 inst_11800 ( .A(net_11059), .Z(net_11648) );
CLKBUF_X2 inst_16039 ( .A(net_15886), .Z(net_15887) );
SDFFR_X2 inst_2565 ( .QN(net_6371), .SE(net_2147), .SI(net_1959), .D(net_778), .CK(net_18129), .RN(x6501) );
CLKBUF_X2 inst_17816 ( .A(net_17663), .Z(net_17664) );
DFFR_X2 inst_7061 ( .QN(net_6328), .D(net_4354), .CK(net_17479), .RN(x6501) );
OAI22_X2 inst_2945 ( .A2(net_4926), .A1(net_2043), .ZN(net_1721), .B2(net_1136), .B1(net_1049) );
SDFF_X2 inst_642 ( .SI(net_8524), .Q(net_8524), .SE(net_3979), .D(net_3965), .CK(net_11085) );
CLKBUF_X2 inst_13035 ( .A(net_12882), .Z(net_12883) );
OAI21_X2 inst_2993 ( .B2(net_5902), .ZN(net_5900), .A(net_5833), .B1(net_698) );
CLKBUF_X2 inst_14736 ( .A(net_14583), .Z(net_14584) );
CLKBUF_X2 inst_13168 ( .A(net_9862), .Z(net_13016) );
SDFF_X2 inst_1018 ( .SI(net_7333), .Q(net_6674), .D(net_6674), .SE(net_3126), .CK(net_11683) );
CLKBUF_X2 inst_18104 ( .A(net_17951), .Z(net_17952) );
CLKBUF_X2 inst_10726 ( .A(net_10573), .Z(net_10574) );
CLKBUF_X2 inst_10655 ( .A(net_9798), .Z(net_10503) );
CLKBUF_X2 inst_16416 ( .A(net_16263), .Z(net_16264) );
CLKBUF_X2 inst_16227 ( .A(net_15002), .Z(net_16075) );
CLKBUF_X2 inst_14160 ( .A(net_9094), .Z(net_14008) );
SDFF_X2 inst_700 ( .Q(net_8433), .D(net_8433), .SI(net_3954), .SE(net_3934), .CK(net_12602) );
CLKBUF_X2 inst_13507 ( .A(net_13354), .Z(net_13355) );
CLKBUF_X2 inst_12295 ( .A(net_10686), .Z(net_12143) );
CLKBUF_X2 inst_13323 ( .A(net_11135), .Z(net_13171) );
AOI22_X2 inst_8107 ( .B1(net_8111), .A1(net_7771), .B2(net_6108), .A2(net_6096), .ZN(net_4040) );
AND2_X2 inst_9152 ( .ZN(net_5589), .A1(net_5588), .A2(net_5462) );
AOI22_X2 inst_8555 ( .ZN(net_2964), .B2(net_2963), .A1(net_2779), .A2(net_2351), .B1(net_903) );
CLKBUF_X2 inst_14457 ( .A(net_14304), .Z(net_14305) );
SDFF_X2 inst_979 ( .SI(net_7314), .Q(net_6721), .D(net_6721), .SE(net_3124), .CK(net_9947) );
NAND2_X2 inst_4568 ( .A2(net_7649), .ZN(net_6082), .A1(net_3081) );
INV_X4 inst_5989 ( .A(net_7436), .ZN(net_3227) );
CLKBUF_X2 inst_9785 ( .A(net_9070), .Z(net_9633) );
SDFFR_X2 inst_2296 ( .SE(net_2260), .Q(net_359), .D(net_359), .CK(net_9321), .RN(x6501), .SI(x1977) );
CLKBUF_X2 inst_13092 ( .A(net_12939), .Z(net_12940) );
CLKBUF_X2 inst_12477 ( .A(net_12324), .Z(net_12325) );
CLKBUF_X2 inst_18883 ( .A(net_13999), .Z(net_18731) );
CLKBUF_X2 inst_17550 ( .A(net_17397), .Z(net_17398) );
CLKBUF_X2 inst_12012 ( .A(net_11859), .Z(net_11860) );
MUX2_X2 inst_4964 ( .A(net_7388), .S(net_2370), .Z(net_2359), .B(net_920) );
CLKBUF_X2 inst_9587 ( .A(net_9434), .Z(net_9435) );
CLKBUF_X2 inst_14133 ( .A(net_13980), .Z(net_13981) );
CLKBUF_X2 inst_14912 ( .A(net_10976), .Z(net_14760) );
CLKBUF_X2 inst_14919 ( .A(net_12298), .Z(net_14767) );
CLKBUF_X2 inst_14802 ( .A(net_14649), .Z(net_14650) );
NAND2_X2 inst_4258 ( .A1(net_7031), .A2(net_5249), .ZN(net_5202) );
AOI22_X2 inst_7889 ( .B1(net_9000), .A2(net_5609), .B2(net_5456), .ZN(net_4542), .A1(net_379) );
CLKBUF_X2 inst_9607 ( .A(net_9454), .Z(net_9455) );
CLKBUF_X2 inst_9764 ( .A(net_9393), .Z(net_9612) );
AOI211_X2 inst_9018 ( .C2(net_2304), .C1(net_2207), .B(net_1925), .ZN(net_1911), .A(net_1910) );
CLKBUF_X2 inst_17537 ( .A(net_17384), .Z(net_17385) );
NAND2_X4 inst_4040 ( .ZN(net_2714), .A2(net_2381), .A1(net_2269) );
SDFF_X2 inst_1059 ( .D(net_7337), .SI(net_6645), .Q(net_6645), .SE(net_3123), .CK(net_9477) );
CLKBUF_X2 inst_18615 ( .A(net_18462), .Z(net_18463) );
CLKBUF_X2 inst_13987 ( .A(net_9848), .Z(net_13835) );
CLKBUF_X2 inst_19117 ( .A(net_15870), .Z(net_18965) );
CLKBUF_X2 inst_16747 ( .A(net_16594), .Z(net_16595) );
CLKBUF_X2 inst_14227 ( .A(net_11276), .Z(net_14075) );
CLKBUF_X2 inst_10215 ( .A(net_10062), .Z(net_10063) );
CLKBUF_X2 inst_16237 ( .A(net_16084), .Z(net_16085) );
NAND2_X2 inst_4328 ( .A1(net_7060), .A2(net_5162), .ZN(net_5129) );
CLKBUF_X2 inst_15240 ( .A(net_13819), .Z(net_15088) );
CLKBUF_X2 inst_15698 ( .A(net_15545), .Z(net_15546) );
NAND2_X2 inst_4173 ( .ZN(net_5336), .A1(net_5083), .A2(net_5082) );
INV_X4 inst_6039 ( .A(net_9014), .ZN(net_1266) );
CLKBUF_X2 inst_17934 ( .A(net_17781), .Z(net_17782) );
CLKBUF_X2 inst_12454 ( .A(net_10187), .Z(net_12302) );
INV_X2 inst_6425 ( .ZN(net_739), .A(net_738) );
SDFF_X2 inst_1104 ( .D(net_7334), .SI(net_6543), .Q(net_6543), .SE(net_3086), .CK(net_12002) );
CLKBUF_X2 inst_17486 ( .A(net_17333), .Z(net_17334) );
SDFFR_X2 inst_2355 ( .SE(net_2757), .D(net_2727), .SI(net_449), .Q(net_449), .CK(net_13849), .RN(x6501) );
CLKBUF_X2 inst_17806 ( .A(net_17653), .Z(net_17654) );
CLKBUF_X2 inst_17756 ( .A(net_17603), .Z(net_17604) );
CLKBUF_X2 inst_10886 ( .A(net_10234), .Z(net_10734) );
INV_X4 inst_5753 ( .A(net_7213), .ZN(net_602) );
DFFR_X2 inst_7058 ( .QN(net_7494), .D(net_4776), .CK(net_17242), .RN(x6501) );
CLKBUF_X2 inst_15794 ( .A(net_15641), .Z(net_15642) );
CLKBUF_X2 inst_12535 ( .A(net_12382), .Z(net_12383) );
CLKBUF_X2 inst_9742 ( .A(net_9589), .Z(net_9590) );
DFFR_X2 inst_7287 ( .QN(net_6344), .D(net_280), .CK(net_16583), .RN(x6501) );
SDFF_X2 inst_574 ( .Q(net_8839), .D(net_8839), .SE(net_3964), .SI(net_3955), .CK(net_10559) );
CLKBUF_X2 inst_12446 ( .A(net_12293), .Z(net_12294) );
CLKBUF_X2 inst_17590 ( .A(net_17437), .Z(net_17438) );
INV_X4 inst_5552 ( .ZN(net_637), .A(x3451) );
CLKBUF_X2 inst_14349 ( .A(net_14196), .Z(net_14197) );
AOI22_X2 inst_8087 ( .B1(net_8040), .A1(net_8006), .B2(net_6102), .A2(net_6097), .ZN(net_4059) );
NAND2_X2 inst_4102 ( .ZN(net_5431), .A2(net_5242), .A1(net_5153) );
SDFF_X2 inst_1229 ( .Q(net_7806), .D(net_7806), .SE(net_2730), .SI(net_2721), .CK(net_15862) );
CLKBUF_X2 inst_10512 ( .A(net_10359), .Z(net_10360) );
CLKBUF_X2 inst_14725 ( .A(net_14572), .Z(net_14573) );
CLKBUF_X2 inst_19031 ( .A(net_18878), .Z(net_18879) );
DFFR_X1 inst_7545 ( .QN(net_5947), .D(net_916), .CK(net_10811), .RN(x6501) );
CLKBUF_X2 inst_13780 ( .A(net_13627), .Z(net_13628) );
CLKBUF_X2 inst_13604 ( .A(net_13451), .Z(net_13452) );
INV_X4 inst_5219 ( .A(net_5783), .ZN(net_5718) );
CLKBUF_X2 inst_18855 ( .A(net_18702), .Z(net_18703) );
CLKBUF_X2 inst_15042 ( .A(net_14889), .Z(net_14890) );
SDFFR_X2 inst_2358 ( .SE(net_2748), .D(net_2725), .SI(net_474), .Q(net_474), .CK(net_16917), .RN(x6501) );
CLKBUF_X2 inst_13139 ( .A(net_12986), .Z(net_12987) );
SDFFR_X2 inst_2125 ( .SI(net_7190), .Q(net_7190), .D(net_6441), .SE(net_4362), .CK(net_17776), .RN(x6501) );
CLKBUF_X2 inst_15827 ( .A(net_15674), .Z(net_15675) );
CLKBUF_X2 inst_17988 ( .A(net_17835), .Z(net_17836) );
CLKBUF_X2 inst_11572 ( .A(net_11419), .Z(net_11420) );
CLKBUF_X2 inst_10549 ( .A(net_10396), .Z(net_10397) );
SDFF_X2 inst_599 ( .SI(net_8392), .Q(net_8392), .SE(net_3969), .D(net_3956), .CK(net_13256) );
CLKBUF_X2 inst_13382 ( .A(net_13229), .Z(net_13230) );
SDFF_X2 inst_541 ( .Q(net_8684), .D(net_8684), .SI(net_3967), .SE(net_3935), .CK(net_10170) );
CLKBUF_X2 inst_16014 ( .A(net_15861), .Z(net_15862) );
NAND2_X4 inst_4047 ( .ZN(net_2508), .A2(net_2222), .A1(net_2088) );
CLKBUF_X2 inst_18645 ( .A(net_18492), .Z(net_18493) );
CLKBUF_X2 inst_13910 ( .A(net_13757), .Z(net_13758) );
SDFF_X2 inst_505 ( .SI(net_8599), .Q(net_8599), .SE(net_3984), .D(net_3947), .CK(net_12460) );
INV_X2 inst_6366 ( .ZN(net_1767), .A(net_1766) );
SDFF_X2 inst_1365 ( .SI(net_7870), .Q(net_7870), .D(net_2704), .SE(net_2558), .CK(net_17017) );
DFFR_X2 inst_7247 ( .QN(net_7307), .D(net_2042), .CK(net_15054), .RN(x6501) );
CLKBUF_X2 inst_15722 ( .A(net_15569), .Z(net_15570) );
AOI22_X2 inst_7936 ( .B1(net_8190), .A1(net_7680), .B2(net_6099), .A2(net_4399), .ZN(net_4188) );
XNOR2_X2 inst_198 ( .ZN(net_1546), .B(net_1183), .A(net_1069) );
CLKBUF_X2 inst_13624 ( .A(net_9820), .Z(net_13472) );
NAND2_X2 inst_4125 ( .ZN(net_5400), .A1(net_5131), .A2(net_5130) );
SDFF_X2 inst_1371 ( .Q(net_8192), .D(net_8192), .SI(net_2574), .SE(net_2561), .CK(net_15603) );
CLKBUF_X2 inst_10809 ( .A(net_10656), .Z(net_10657) );
INV_X4 inst_5622 ( .A(net_8956), .ZN(net_1450) );
NAND2_X2 inst_4321 ( .A1(net_7099), .A2(net_5164), .ZN(net_5136) );
SDFF_X2 inst_1644 ( .SI(net_7720), .Q(net_7720), .D(net_2575), .SE(net_2559), .CK(net_15986) );
INV_X2 inst_6346 ( .ZN(net_2421), .A(net_2353) );
CLKBUF_X2 inst_18531 ( .A(net_15667), .Z(net_18379) );
CLKBUF_X2 inst_12645 ( .A(net_12492), .Z(net_12493) );
CLKBUF_X2 inst_18921 ( .A(net_18768), .Z(net_18769) );
AOI21_X2 inst_8946 ( .B2(net_5871), .ZN(net_5601), .A(net_5600), .B1(x521) );
DFFR_X1 inst_7529 ( .Q(net_7659), .D(net_7655), .CK(net_12715), .RN(x6501) );
CLKBUF_X2 inst_13333 ( .A(net_13180), .Z(net_13181) );
CLKBUF_X2 inst_9351 ( .A(net_9113), .Z(net_9199) );
CLKBUF_X2 inst_16194 ( .A(net_11998), .Z(net_16042) );
CLKBUF_X2 inst_15071 ( .A(net_14918), .Z(net_14919) );
CLKBUF_X2 inst_17335 ( .A(net_17182), .Z(net_17183) );
NOR2_X2 inst_3511 ( .ZN(net_2007), .A2(net_1820), .A1(net_1535) );
CLKBUF_X2 inst_18168 ( .A(net_10653), .Z(net_18016) );
DFF_X1 inst_6726 ( .Q(net_6772), .D(net_5643), .CK(net_9257) );
CLKBUF_X2 inst_10363 ( .A(net_9847), .Z(net_10211) );
INV_X4 inst_5693 ( .A(net_5959), .ZN(x2746) );
CLKBUF_X2 inst_9992 ( .A(net_9839), .Z(net_9840) );
XNOR2_X2 inst_263 ( .B(net_8891), .ZN(net_1157), .A(net_1156) );
CLKBUF_X2 inst_18352 ( .A(net_17306), .Z(net_18200) );
CLKBUF_X2 inst_10889 ( .A(net_10736), .Z(net_10737) );
CLKBUF_X2 inst_15831 ( .A(net_15678), .Z(net_15679) );
DFFR_X1 inst_7399 ( .D(net_5757), .CK(net_16771), .RN(x6501), .Q(x494) );
INV_X4 inst_5953 ( .A(net_8905), .ZN(net_2790) );
DFF_X1 inst_6742 ( .Q(net_6786), .D(net_5627), .CK(net_11420) );
INV_X2 inst_6307 ( .ZN(net_3897), .A(net_3594) );
DFFR_X1 inst_7371 ( .QN(net_6313), .D(net_5883), .CK(net_14066), .RN(x6501) );
CLKBUF_X2 inst_10650 ( .A(net_10131), .Z(net_10498) );
CLKBUF_X2 inst_10121 ( .A(net_9968), .Z(net_9969) );
CLKBUF_X2 inst_11923 ( .A(net_11621), .Z(net_11771) );
NAND2_X2 inst_4118 ( .ZN(net_5409), .A1(net_5231), .A2(net_5008) );
CLKBUF_X2 inst_13410 ( .A(net_13257), .Z(net_13258) );
INV_X4 inst_5440 ( .ZN(net_1090), .A(net_865) );
NAND2_X2 inst_4849 ( .A1(net_8279), .ZN(net_901), .A2(net_562) );
CLKBUF_X2 inst_14689 ( .A(net_14536), .Z(net_14537) );
CLKBUF_X2 inst_17504 ( .A(net_17351), .Z(net_17352) );
CLKBUF_X2 inst_16593 ( .A(net_16440), .Z(net_16441) );
AOI22_X2 inst_8185 ( .B1(net_8568), .A1(net_8457), .A2(net_6263), .B2(net_6262), .ZN(net_3847) );
CLKBUF_X2 inst_11223 ( .A(net_11070), .Z(net_11071) );
CLKBUF_X2 inst_17647 ( .A(net_17494), .Z(net_17495) );
DFFR_X1 inst_7413 ( .QN(net_6342), .D(net_5737), .CK(net_14226), .RN(x6501) );
CLKBUF_X2 inst_15709 ( .A(net_15556), .Z(net_15557) );
CLKBUF_X2 inst_14263 ( .A(net_11202), .Z(net_14111) );
AOI222_X1 inst_8698 ( .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3053), .B1(net_3052), .C1(net_3051), .A2(net_2871) );
INV_X8 inst_5034 ( .ZN(net_1561), .A(net_836) );
NAND2_X2 inst_4853 ( .A2(net_7410), .A1(net_1236), .ZN(net_893) );
INV_X2 inst_6322 ( .ZN(net_3341), .A(net_3285) );
NAND3_X2 inst_3898 ( .ZN(net_5640), .A1(net_5569), .A3(net_5503), .A2(net_5402) );
CLKBUF_X2 inst_17083 ( .A(net_16930), .Z(net_16931) );
INV_X4 inst_5254 ( .A(net_2450), .ZN(net_2333) );
CLKBUF_X2 inst_18569 ( .A(net_18416), .Z(net_18417) );
CLKBUF_X2 inst_18161 ( .A(net_10115), .Z(net_18009) );
CLKBUF_X2 inst_9370 ( .A(net_9217), .Z(net_9218) );
CLKBUF_X2 inst_11949 ( .A(net_11067), .Z(net_11797) );
NOR2_X2 inst_3503 ( .A2(net_2397), .ZN(net_2342), .A1(net_1862) );
CLKBUF_X2 inst_13974 ( .A(net_13821), .Z(net_13822) );
CLKBUF_X2 inst_15836 ( .A(net_15683), .Z(net_15684) );
AOI22_X2 inst_7973 ( .B1(net_8162), .A1(net_7720), .B2(net_6101), .A2(net_6095), .ZN(net_6006) );
NAND2_X2 inst_4138 ( .ZN(net_5383), .A2(net_5218), .A1(net_5117) );
XOR2_X2 inst_52 ( .A(net_3274), .Z(net_996), .B(net_594) );
CLKBUF_X2 inst_12600 ( .A(net_12447), .Z(net_12448) );
SDFF_X2 inst_668 ( .Q(net_8443), .D(net_8443), .SI(net_3949), .SE(net_3934), .CK(net_12609) );
CLKBUF_X2 inst_17799 ( .A(net_17646), .Z(net_17647) );
OAI21_X2 inst_3049 ( .B2(net_8230), .B1(net_4850), .ZN(net_4762), .A(net_2615) );
CLKBUF_X2 inst_15804 ( .A(net_14763), .Z(net_15652) );
CLKBUF_X2 inst_11987 ( .A(net_11834), .Z(net_11835) );
CLKBUF_X2 inst_16015 ( .A(net_12179), .Z(net_15863) );
CLKBUF_X2 inst_17571 ( .A(net_9497), .Z(net_17419) );
NAND2_X2 inst_4159 ( .ZN(net_5355), .A1(net_5098), .A2(net_5097) );
CLKBUF_X2 inst_12567 ( .A(net_10885), .Z(net_12415) );
NOR2_X2 inst_3349 ( .ZN(net_5576), .A1(net_5432), .A2(net_5431) );
CLKBUF_X2 inst_11444 ( .A(net_9556), .Z(net_11292) );
CLKBUF_X2 inst_10057 ( .A(net_9904), .Z(net_9905) );
SDFFR_X2 inst_2545 ( .QN(net_6349), .SE(net_2147), .SI(net_1612), .D(net_970), .CK(net_14955), .RN(x6501) );
AOI22_X2 inst_8220 ( .B1(net_8573), .A1(net_8462), .A2(net_6263), .B2(net_6262), .ZN(net_3816) );
CLKBUF_X2 inst_18441 ( .A(net_18288), .Z(net_18289) );
CLKBUF_X2 inst_12390 ( .A(net_10708), .Z(net_12238) );
CLKBUF_X2 inst_10722 ( .A(net_10569), .Z(net_10570) );
AOI22_X2 inst_7999 ( .B1(net_8029), .A1(net_7995), .B2(net_6102), .A2(net_6097), .ZN(net_4134) );
CLKBUF_X2 inst_13077 ( .A(net_12924), .Z(net_12925) );
SDFFR_X1 inst_2768 ( .Q(net_7296), .SI(net_7260), .D(net_2129), .SE(net_1327), .CK(net_18249), .RN(x6501) );
CLKBUF_X2 inst_14657 ( .A(net_14504), .Z(net_14505) );
CLKBUF_X2 inst_17459 ( .A(net_17306), .Z(net_17307) );
CLKBUF_X2 inst_9878 ( .A(net_9725), .Z(net_9726) );
SDFF_X2 inst_1835 ( .D(net_7263), .SI(net_6880), .Q(net_6880), .SE(net_6284), .CK(net_14348) );
CLKBUF_X2 inst_16890 ( .A(net_11003), .Z(net_16738) );
CLKBUF_X2 inst_19183 ( .A(net_13526), .Z(net_19031) );
CLKBUF_X2 inst_15861 ( .A(net_15708), .Z(net_15709) );
CLKBUF_X2 inst_13777 ( .A(net_13624), .Z(net_13625) );
CLKBUF_X2 inst_15614 ( .A(net_15461), .Z(net_15462) );
NAND2_X2 inst_4639 ( .ZN(net_2441), .A2(net_2440), .A1(net_2346) );
CLKBUF_X2 inst_12399 ( .A(net_11636), .Z(net_12247) );
CLKBUF_X2 inst_9670 ( .A(net_9517), .Z(net_9518) );
AOI22_X2 inst_7797 ( .B1(net_7186), .A2(net_6129), .B2(net_5655), .ZN(net_4792), .A1(net_1296) );
CLKBUF_X2 inst_15410 ( .A(net_15257), .Z(net_15258) );
CLKBUF_X2 inst_15176 ( .A(net_15023), .Z(net_15024) );
SDFF_X2 inst_621 ( .SI(net_8532), .Q(net_8532), .SE(net_3979), .D(net_3966), .CK(net_10926) );
AOI22_X2 inst_7764 ( .B1(net_6991), .A1(net_6951), .A2(net_5443), .B2(net_5442), .ZN(net_5350) );
CLKBUF_X2 inst_18386 ( .A(net_18233), .Z(net_18234) );
SDFFR_X2 inst_2560 ( .Q(net_6386), .D(net_6386), .SE(net_2147), .SI(net_1461), .CK(net_18234), .RN(x6501) );
CLKBUF_X2 inst_17188 ( .A(net_17035), .Z(net_17036) );
CLKBUF_X2 inst_15224 ( .A(net_15071), .Z(net_15072) );
CLKBUF_X2 inst_12236 ( .A(net_12083), .Z(net_12084) );
CLKBUF_X2 inst_9651 ( .A(net_9498), .Z(net_9499) );
CLKBUF_X2 inst_14435 ( .A(net_14282), .Z(net_14283) );
SDFF_X2 inst_1387 ( .SI(net_7291), .Q(net_7108), .D(net_7108), .SE(net_6278), .CK(net_17716) );
CLKBUF_X2 inst_15138 ( .A(net_9380), .Z(net_14986) );
CLKBUF_X2 inst_13687 ( .A(net_12558), .Z(net_13535) );
SDFFR_X2 inst_2365 ( .SE(net_2260), .Q(net_333), .D(net_333), .CK(net_9305), .RN(x6501), .SI(x2494) );
CLKBUF_X2 inst_18367 ( .A(net_18214), .Z(net_18215) );
CLKBUF_X2 inst_16851 ( .A(net_16698), .Z(net_16699) );
CLKBUF_X2 inst_12094 ( .A(net_11941), .Z(net_11942) );
SDFFR_X2 inst_2250 ( .D(net_7396), .SE(net_2801), .SI(net_205), .Q(net_205), .CK(net_14768), .RN(x6501) );
CLKBUF_X2 inst_15190 ( .A(net_14146), .Z(net_15038) );
INV_X16 inst_6629 ( .ZN(net_3857), .A(net_3380) );
SDFFR_X2 inst_2187 ( .QN(net_7411), .SE(net_2778), .SI(net_2777), .D(net_2021), .CK(net_17947), .RN(x6501) );
CLKBUF_X2 inst_13221 ( .A(net_13068), .Z(net_13069) );
CLKBUF_X2 inst_11215 ( .A(net_10278), .Z(net_11063) );
INV_X4 inst_5747 ( .A(net_6390), .ZN(net_1308) );
CLKBUF_X2 inst_14323 ( .A(net_14170), .Z(net_14171) );
DFFR_X1 inst_7448 ( .QN(net_8931), .D(net_4751), .CK(net_14851), .RN(x6501) );
XOR2_X2 inst_25 ( .A(net_1776), .Z(net_1360), .B(net_830) );
AND3_X4 inst_9043 ( .ZN(net_2440), .A1(net_2278), .A3(net_1976), .A2(net_1596) );
INV_X4 inst_5239 ( .A(net_2489), .ZN(net_2014) );
INV_X8 inst_5032 ( .ZN(net_2453), .A(net_2210) );
INV_X4 inst_5166 ( .ZN(net_6175), .A(net_3081) );
CLKBUF_X2 inst_16210 ( .A(net_16057), .Z(net_16058) );
CLKBUF_X2 inst_9691 ( .A(net_9538), .Z(net_9539) );
SDFFR_X2 inst_2500 ( .Q(net_8993), .D(net_8993), .SI(net_4551), .SE(net_2562), .CK(net_17266), .RN(x6501) );
CLKBUF_X2 inst_12119 ( .A(net_10804), .Z(net_11967) );
CLKBUF_X2 inst_9734 ( .A(net_9581), .Z(net_9582) );
NAND2_X2 inst_4395 ( .A1(net_7125), .A2(net_5166), .ZN(net_5062) );
NOR2_X2 inst_3434 ( .A2(net_3093), .ZN(net_3075), .A1(net_1850) );
NAND2_X2 inst_4296 ( .A1(net_7131), .A2(net_5166), .ZN(net_5161) );
OAI211_X2 inst_3204 ( .C2(net_7222), .ZN(net_2399), .B(net_2085), .A(net_2084), .C1(net_2074) );
CLKBUF_X2 inst_14219 ( .A(net_9150), .Z(net_14067) );
NOR2_X2 inst_3421 ( .ZN(net_3216), .A1(net_3176), .A2(net_3157) );
NAND2_X2 inst_4444 ( .A1(net_6844), .A2(net_5016), .ZN(net_4983) );
CLKBUF_X2 inst_12019 ( .A(net_11866), .Z(net_11867) );
SDFFR_X1 inst_2679 ( .SI(net_7543), .SE(net_5043), .CK(net_9704), .RN(x6501), .Q(x4023), .D(x4023) );
DFFS_X1 inst_6935 ( .D(net_6145), .CK(net_13657), .SN(x6501), .Q(x697) );
NAND3_X2 inst_3949 ( .A3(net_6207), .ZN(net_4393), .A1(net_4323), .A2(net_4322) );
CLKBUF_X2 inst_15731 ( .A(net_15578), .Z(net_15579) );
CLKBUF_X2 inst_16727 ( .A(net_12217), .Z(net_16575) );
NAND2_X2 inst_4617 ( .A2(net_6144), .ZN(net_2607), .A1(net_2606) );
SDFF_X2 inst_1777 ( .D(net_7282), .SI(net_6859), .Q(net_6859), .SE(net_6282), .CK(net_14898) );
CLKBUF_X2 inst_18919 ( .A(net_18766), .Z(net_18767) );
CLKBUF_X2 inst_14971 ( .A(net_14818), .Z(net_14819) );
SDFF_X2 inst_1068 ( .D(net_7329), .SI(net_6538), .Q(net_6538), .SE(net_3086), .CK(net_11285) );
SDFF_X2 inst_886 ( .Q(net_8565), .D(net_8565), .SI(net_3946), .SE(net_3878), .CK(net_11042) );
CLKBUF_X2 inst_12799 ( .A(net_12646), .Z(net_12647) );
CLKBUF_X2 inst_11799 ( .A(net_10828), .Z(net_11647) );
CLKBUF_X2 inst_16608 ( .A(net_16455), .Z(net_16456) );
CLKBUF_X2 inst_12509 ( .A(net_12207), .Z(net_12357) );
CLKBUF_X2 inst_15409 ( .A(net_15256), .Z(net_15257) );
INV_X4 inst_5350 ( .ZN(net_4926), .A(net_4924) );
CLKBUF_X2 inst_18620 ( .A(net_18467), .Z(net_18468) );
CLKBUF_X2 inst_15251 ( .A(net_15098), .Z(net_15099) );
CLKBUF_X2 inst_13319 ( .A(net_13166), .Z(net_13167) );
NAND2_X2 inst_4468 ( .ZN(net_4727), .A2(net_4725), .A1(net_4505) );
CLKBUF_X2 inst_11740 ( .A(net_11587), .Z(net_11588) );
CLKBUF_X2 inst_11533 ( .A(net_11380), .Z(net_11381) );
CLKBUF_X2 inst_14450 ( .A(net_11116), .Z(net_14298) );
CLKBUF_X2 inst_11484 ( .A(net_10040), .Z(net_11332) );
CLKBUF_X2 inst_17520 ( .A(net_10580), .Z(net_17368) );
CLKBUF_X2 inst_11270 ( .A(net_10368), .Z(net_11118) );
CLKBUF_X2 inst_15874 ( .A(net_15721), .Z(net_15722) );
CLKBUF_X2 inst_12380 ( .A(net_11141), .Z(net_12228) );
AOI221_X2 inst_8844 ( .C1(net_8154), .B1(net_7712), .C2(net_6101), .B2(net_6095), .ZN(net_6060), .A(net_4278) );
SDFF_X2 inst_1969 ( .D(net_7265), .SI(net_6882), .Q(net_6882), .SE(net_6284), .CK(net_14314) );
AOI22_X2 inst_7837 ( .A2(net_6453), .A1(net_5654), .B2(net_5595), .ZN(net_4674), .B1(net_335) );
CLKBUF_X2 inst_11382 ( .A(net_10879), .Z(net_11230) );
AND2_X4 inst_9128 ( .ZN(net_1391), .A2(net_889), .A1(net_164) );
CLKBUF_X2 inst_15631 ( .A(net_15478), .Z(net_15479) );
CLKBUF_X2 inst_9348 ( .A(net_9195), .Z(net_9196) );
AOI22_X2 inst_8183 ( .A1(net_8605), .B1(net_8420), .A2(net_3864), .B2(net_3863), .ZN(net_3849) );
DFFS_X1 inst_6914 ( .Q(net_6335), .D(net_5725), .CK(net_14211), .SN(x6501) );
CLKBUF_X2 inst_15004 ( .A(net_14229), .Z(net_14852) );
CLKBUF_X2 inst_18993 ( .A(net_18840), .Z(net_18841) );
INV_X2 inst_6540 ( .A(net_6356), .ZN(net_2121) );
CLKBUF_X2 inst_14536 ( .A(net_14383), .Z(net_14384) );
CLKBUF_X2 inst_18928 ( .A(net_14072), .Z(net_18776) );
CLKBUF_X2 inst_13136 ( .A(net_9060), .Z(net_12984) );
OAI21_X2 inst_3150 ( .ZN(net_1986), .A(net_1985), .B2(net_1984), .B1(net_721) );
CLKBUF_X2 inst_10761 ( .A(net_10608), .Z(net_10609) );
CLKBUF_X2 inst_18793 ( .A(net_14949), .Z(net_18641) );
CLKBUF_X2 inst_15976 ( .A(net_12847), .Z(net_15824) );
CLKBUF_X2 inst_12765 ( .A(net_12612), .Z(net_12613) );
AOI22_X2 inst_8522 ( .B1(net_6655), .A1(net_6622), .A2(net_6213), .B2(net_6138), .ZN(net_3418) );
CLKBUF_X2 inst_14741 ( .A(net_14588), .Z(net_14589) );
INV_X2 inst_6216 ( .ZN(net_5494), .A(net_5365) );
INV_X4 inst_5791 ( .A(net_9006), .ZN(net_2656) );
SDFF_X2 inst_866 ( .Q(net_8557), .D(net_8557), .SI(net_3943), .SE(net_3878), .CK(net_13307) );
CLKBUF_X2 inst_11061 ( .A(net_10908), .Z(net_10909) );
SDFF_X2 inst_1439 ( .SI(net_7264), .Q(net_7081), .D(net_7081), .SE(net_6278), .CK(net_14366) );
DFFR_X2 inst_7214 ( .D(net_2355), .QN(net_228), .CK(net_18175), .RN(x6501) );
NAND4_X2 inst_3640 ( .ZN(net_5021), .A2(net_4807), .A4(net_4706), .A3(net_4645), .A1(net_4478) );
CLKBUF_X2 inst_12367 ( .A(net_12214), .Z(net_12215) );
AOI22_X2 inst_8444 ( .B1(net_6535), .A1(net_6502), .A2(net_6137), .B2(net_6104), .ZN(net_3497) );
CLKBUF_X2 inst_17950 ( .A(net_17797), .Z(net_17798) );
CLKBUF_X2 inst_17200 ( .A(net_17047), .Z(net_17048) );
INV_X4 inst_5604 ( .A(net_7385), .ZN(net_972) );
XNOR2_X2 inst_248 ( .ZN(net_1203), .A(net_1202), .B(net_490) );
OAI21_X2 inst_3107 ( .ZN(net_2490), .B2(net_2489), .A(net_2330), .B1(net_1847) );
SDFF_X2 inst_1919 ( .SI(net_7036), .Q(net_7036), .SE(net_6277), .D(net_2544), .CK(net_15869) );
CLKBUF_X2 inst_15747 ( .A(net_14156), .Z(net_15595) );
CLKBUF_X2 inst_18442 ( .A(net_18289), .Z(net_18290) );
CLKBUF_X2 inst_12222 ( .A(net_12069), .Z(net_12070) );
CLKBUF_X2 inst_18238 ( .A(net_18085), .Z(net_18086) );
CLKBUF_X2 inst_10528 ( .A(net_10375), .Z(net_10376) );
CLKBUF_X2 inst_15938 ( .A(net_15785), .Z(net_15786) );
CLKBUF_X2 inst_18508 ( .A(net_18355), .Z(net_18356) );
SDFF_X2 inst_1960 ( .D(net_7267), .SI(net_6964), .Q(net_6964), .SE(net_6283), .CK(net_14075) );
CLKBUF_X2 inst_15675 ( .A(net_15522), .Z(net_15523) );
AOI221_X4 inst_8712 ( .C1(net_8182), .B1(net_7672), .C2(net_6099), .ZN(net_6047), .B2(net_4399), .A(net_4288) );
CLKBUF_X2 inst_13273 ( .A(net_13120), .Z(net_13121) );
CLKBUF_X2 inst_11886 ( .A(net_9450), .Z(net_11734) );
CLKBUF_X2 inst_10283 ( .A(net_10130), .Z(net_10131) );
CLKBUF_X2 inst_10659 ( .A(net_10506), .Z(net_10507) );
CLKBUF_X2 inst_10744 ( .A(net_10591), .Z(net_10592) );
NAND2_X2 inst_4636 ( .ZN(net_2577), .A2(net_2260), .A1(net_2091) );
XNOR2_X2 inst_302 ( .ZN(net_977), .A(net_976), .B(net_975) );
SDFF_X2 inst_673 ( .Q(net_8412), .D(net_8412), .SI(net_3938), .SE(net_3934), .CK(net_13039) );
NOR2_X2 inst_3585 ( .A2(net_7221), .ZN(net_1619), .A1(net_584) );
SDFF_X2 inst_1151 ( .SI(net_7332), .Q(net_6607), .D(net_6607), .SE(net_3069), .CK(net_9412) );
CLKBUF_X2 inst_14952 ( .A(net_14799), .Z(net_14800) );
CLKBUF_X2 inst_11399 ( .A(net_10590), .Z(net_11247) );
SDFF_X2 inst_561 ( .Q(net_8676), .D(net_8676), .SI(net_3946), .SE(net_3935), .CK(net_11089) );
CLKBUF_X2 inst_13417 ( .A(net_13264), .Z(net_13265) );
CLKBUF_X2 inst_12999 ( .A(net_10294), .Z(net_12847) );
CLKBUF_X2 inst_10903 ( .A(net_10453), .Z(net_10751) );
SDFFR_X2 inst_2505 ( .Q(net_8976), .D(net_8976), .SI(net_2622), .SE(net_2562), .CK(net_16625), .RN(x6501) );
INV_X2 inst_6504 ( .A(net_7422), .ZN(net_539) );
CLKBUF_X2 inst_12253 ( .A(net_12100), .Z(net_12101) );
SDFF_X2 inst_1641 ( .SI(net_7715), .Q(net_7715), .D(net_2706), .SE(net_2559), .CK(net_18852) );
DFF_X1 inst_6765 ( .Q(net_7545), .D(net_4607), .CK(net_9723) );
CLKBUF_X2 inst_19167 ( .A(net_19014), .Z(net_19015) );
CLKBUF_X2 inst_12524 ( .A(net_12371), .Z(net_12372) );
CLKBUF_X2 inst_14620 ( .A(net_12793), .Z(net_14468) );
CLKBUF_X2 inst_11749 ( .A(net_9915), .Z(net_11597) );
XNOR2_X2 inst_196 ( .ZN(net_1548), .B(net_1196), .A(net_1184) );
SDFF_X2 inst_1567 ( .Q(net_8129), .D(net_8129), .SI(net_2719), .SE(net_2541), .CK(net_18789) );
CLKBUF_X2 inst_18661 ( .A(net_18508), .Z(net_18509) );
CLKBUF_X2 inst_17542 ( .A(net_10743), .Z(net_17390) );
CLKBUF_X2 inst_15161 ( .A(net_11632), .Z(net_15009) );
NOR2_X2 inst_3451 ( .ZN(net_2939), .A2(net_2838), .A1(net_1800) );
SDFFR_X2 inst_2417 ( .D(net_2687), .SE(net_2313), .SI(net_462), .Q(net_462), .CK(net_16915), .RN(x6501) );
CLKBUF_X2 inst_13481 ( .A(net_12213), .Z(net_13329) );
CLKBUF_X2 inst_12828 ( .A(net_12493), .Z(net_12676) );
AOI22_X2 inst_8405 ( .A1(net_8601), .B1(net_8416), .A2(net_3864), .B2(net_3863), .ZN(net_3647) );
CLKBUF_X2 inst_17960 ( .A(net_13810), .Z(net_17808) );
INV_X4 inst_5606 ( .A(net_7424), .ZN(net_3194) );
CLKBUF_X2 inst_14371 ( .A(net_14218), .Z(net_14219) );
XNOR2_X2 inst_298 ( .B(net_1226), .ZN(net_984), .A(net_507) );
SDFFR_X2 inst_2180 ( .QN(net_7586), .D(net_3954), .SE(net_3144), .SI(net_491), .CK(net_12648), .RN(x6501) );
SDFF_X2 inst_1856 ( .D(net_7283), .SI(net_6940), .Q(net_6940), .SE(net_6281), .CK(net_18988) );
CLKBUF_X2 inst_9379 ( .A(net_9087), .Z(net_9227) );
INV_X4 inst_5507 ( .A(net_908), .ZN(net_857) );
CLKBUF_X2 inst_15993 ( .A(net_15840), .Z(net_15841) );
INV_X2 inst_6594 ( .A(net_6127), .ZN(net_6126) );
CLKBUF_X2 inst_11390 ( .A(net_11237), .Z(net_11238) );
CLKBUF_X2 inst_11124 ( .A(net_9912), .Z(net_10972) );
INV_X2 inst_6180 ( .ZN(net_5870), .A(net_5825) );
NOR2_X2 inst_3529 ( .ZN(net_1713), .A2(net_1636), .A1(net_701) );
CLKBUF_X2 inst_14548 ( .A(net_12430), .Z(net_14396) );
SDFF_X2 inst_2040 ( .SI(net_7788), .Q(net_7788), .D(net_2575), .SE(net_2459), .CK(net_15945) );
CLKBUF_X2 inst_10834 ( .A(net_10681), .Z(net_10682) );
CLKBUF_X2 inst_17956 ( .A(net_17803), .Z(net_17804) );
DFFR_X2 inst_7327 ( .QN(net_6806), .D(net_6803), .CK(net_9635), .RN(x6501) );
NAND2_X2 inst_4742 ( .ZN(net_2718), .A2(net_1586), .A1(net_1144) );
CLKBUF_X2 inst_18820 ( .A(net_10091), .Z(net_18668) );
INV_X2 inst_6527 ( .A(net_6358), .ZN(net_2132) );
INV_X4 inst_6099 ( .A(net_6477), .ZN(net_911) );
CLKBUF_X2 inst_12687 ( .A(net_12534), .Z(net_12535) );
NAND2_X2 inst_4561 ( .ZN(net_3230), .A1(net_3187), .A2(net_3152) );
CLKBUF_X2 inst_11315 ( .A(net_11162), .Z(net_11163) );
CLKBUF_X2 inst_9324 ( .A(net_9112), .Z(net_9172) );
CLKBUF_X2 inst_9611 ( .A(net_9344), .Z(net_9459) );
INV_X2 inst_6221 ( .ZN(net_5489), .A(net_5345) );
SDFFR_X1 inst_2743 ( .SI(net_9022), .Q(net_9022), .D(net_7451), .SE(net_3208), .CK(net_12834), .RN(x6501) );
CLKBUF_X2 inst_17978 ( .A(net_17825), .Z(net_17826) );
SDFFS_X2 inst_2083 ( .SI(net_7376), .SE(net_2794), .Q(net_165), .D(net_165), .CK(net_17728), .SN(x6501) );
CLKBUF_X2 inst_15144 ( .A(net_14991), .Z(net_14992) );
SDFF_X2 inst_1470 ( .SI(net_7295), .Q(net_7152), .D(net_7152), .SE(net_6279), .CK(net_18199) );
CLKBUF_X2 inst_17493 ( .A(net_10249), .Z(net_17341) );
AOI22_X2 inst_8019 ( .B1(net_7929), .A1(net_7827), .B2(net_6103), .A2(net_4398), .ZN(net_4117) );
CLKBUF_X2 inst_16198 ( .A(net_16045), .Z(net_16046) );
CLKBUF_X2 inst_16294 ( .A(net_11591), .Z(net_16142) );
SDFF_X2 inst_1213 ( .Q(net_7967), .D(net_7967), .SE(net_2755), .SI(net_2711), .CK(net_14303) );
OAI21_X2 inst_3072 ( .ZN(net_4224), .A(net_4222), .B2(net_4221), .B1(net_732) );
DFFR_X1 inst_7524 ( .D(net_1294), .Q(net_299), .CK(net_16604), .RN(x6501) );
CLKBUF_X2 inst_12128 ( .A(net_10991), .Z(net_11976) );
CLKBUF_X2 inst_14094 ( .A(net_13941), .Z(net_13942) );
SDFFR_X2 inst_2452 ( .D(net_7511), .SE(net_2313), .SI(net_427), .Q(net_427), .CK(net_14546), .RN(x6501) );
CLKBUF_X2 inst_11370 ( .A(net_10371), .Z(net_11218) );
CLKBUF_X2 inst_17243 ( .A(net_17090), .Z(net_17091) );
SDFF_X2 inst_428 ( .Q(net_8755), .D(net_8755), .SE(net_3982), .SI(net_3959), .CK(net_10194) );
CLKBUF_X2 inst_11821 ( .A(net_11668), .Z(net_11669) );
CLKBUF_X2 inst_17842 ( .A(net_17689), .Z(net_17690) );
AND2_X4 inst_9093 ( .ZN(net_2730), .A2(net_2381), .A1(net_2261) );
CLKBUF_X2 inst_17043 ( .A(net_10720), .Z(net_16891) );
XOR2_X1 inst_97 ( .Z(net_1386), .B(net_1385), .A(net_708) );
CLKBUF_X2 inst_15658 ( .A(net_15505), .Z(net_15506) );
SDFF_X2 inst_775 ( .Q(net_8787), .D(net_8787), .SI(net_3946), .SE(net_3879), .CK(net_11051) );
AOI22_X2 inst_8120 ( .A1(net_7946), .B1(net_7776), .A2(net_6092), .B2(net_6091), .ZN(net_4029) );
NAND2_X2 inst_4652 ( .ZN(net_2297), .A1(net_2296), .A2(net_2212) );
CLKBUF_X2 inst_16058 ( .A(net_15905), .Z(net_15906) );
CLKBUF_X2 inst_18815 ( .A(net_18662), .Z(net_18663) );
CLKBUF_X2 inst_18446 ( .A(net_18293), .Z(net_18294) );
CLKBUF_X2 inst_11102 ( .A(net_10949), .Z(net_10950) );
CLKBUF_X2 inst_11812 ( .A(net_11440), .Z(net_11660) );
CLKBUF_X2 inst_14281 ( .A(net_12053), .Z(net_14129) );
CLKBUF_X2 inst_17020 ( .A(net_16867), .Z(net_16868) );
CLKBUF_X2 inst_15124 ( .A(net_14971), .Z(net_14972) );
SDFFR_X2 inst_2242 ( .Q(net_7457), .D(net_7457), .SE(net_2863), .CK(net_10615), .SI(x13527), .RN(x6501) );
CLKBUF_X2 inst_12954 ( .A(net_10983), .Z(net_12802) );
SDFF_X2 inst_1671 ( .SI(net_7770), .Q(net_7770), .D(net_2656), .SE(net_2560), .CK(net_14399) );
NAND2_X2 inst_4581 ( .A2(net_4362), .ZN(net_2954), .A1(net_2953) );
CLKBUF_X2 inst_10044 ( .A(net_9891), .Z(net_9892) );
CLKBUF_X2 inst_13203 ( .A(net_13050), .Z(net_13051) );
OR2_X2 inst_2884 ( .A1(net_2244), .ZN(net_1822), .A2(net_1821) );
SDFF_X2 inst_600 ( .SI(net_8393), .Q(net_8393), .SE(net_3969), .D(net_3963), .CK(net_10933) );
CLKBUF_X2 inst_13662 ( .A(net_13509), .Z(net_13510) );
CLKBUF_X2 inst_15906 ( .A(net_14606), .Z(net_15754) );
INV_X4 inst_5319 ( .ZN(net_4404), .A(net_1432) );
NAND2_X2 inst_4498 ( .ZN(net_4472), .A2(net_4468), .A1(net_4404) );
SDFF_X2 inst_1194 ( .D(net_7319), .SI(net_6528), .Q(net_6528), .SE(net_3086), .CK(net_9826) );
CLKBUF_X2 inst_14292 ( .A(net_14139), .Z(net_14140) );
XOR2_X2 inst_49 ( .B(net_3113), .Z(net_1012), .A(net_1011) );
CLKBUF_X2 inst_14353 ( .A(net_14200), .Z(net_14201) );
CLKBUF_X2 inst_17196 ( .A(net_17043), .Z(net_17044) );
CLKBUF_X2 inst_14288 ( .A(net_14135), .Z(net_14136) );
CLKBUF_X2 inst_15306 ( .A(net_11779), .Z(net_15154) );
NAND2_X2 inst_4097 ( .ZN(net_5437), .A1(net_5245), .A2(net_5015) );
SDFF_X2 inst_693 ( .Q(net_8875), .D(net_8875), .SI(net_3942), .SE(net_3936), .CK(net_10538) );
CLKBUF_X2 inst_18439 ( .A(net_12499), .Z(net_18287) );
CLKBUF_X2 inst_17246 ( .A(net_16157), .Z(net_17094) );
CLKBUF_X2 inst_10119 ( .A(net_9966), .Z(net_9967) );
AOI21_X2 inst_8920 ( .B2(net_5843), .ZN(net_5716), .A(net_5715), .B1(x258) );
INV_X2 inst_6217 ( .ZN(net_5493), .A(net_5361) );
DFFR_X1 inst_7383 ( .D(net_5877), .CK(net_17183), .RN(x6501), .Q(x225) );
DFFR_X1 inst_7390 ( .D(net_5859), .CK(net_16781), .RN(x6501), .Q(x434) );
CLKBUF_X2 inst_17402 ( .A(net_17249), .Z(net_17250) );
AOI22_X2 inst_8303 ( .B1(net_8843), .A1(net_8362), .A2(net_6265), .B2(net_6253), .ZN(net_6068) );
CLKBUF_X2 inst_18605 ( .A(net_15969), .Z(net_18453) );
CLKBUF_X2 inst_14987 ( .A(net_14834), .Z(net_14835) );
SDFF_X2 inst_908 ( .SI(net_8726), .Q(net_8726), .SE(net_6195), .D(net_3963), .CK(net_10888) );
CLKBUF_X2 inst_11690 ( .A(net_11537), .Z(net_11538) );
CLKBUF_X2 inst_13731 ( .A(net_13578), .Z(net_13579) );
CLKBUF_X2 inst_9227 ( .A(net_9074), .Z(net_9075) );
XNOR2_X2 inst_218 ( .B(net_8891), .ZN(net_1408), .A(net_1407) );
NAND4_X2 inst_3647 ( .ZN(net_4914), .A3(net_4653), .A2(net_4523), .A4(net_4521), .A1(net_4460) );
CLKBUF_X2 inst_14773 ( .A(net_14620), .Z(net_14621) );
CLKBUF_X2 inst_11865 ( .A(net_9565), .Z(net_11713) );
CLKBUF_X2 inst_18094 ( .A(net_17941), .Z(net_17942) );
CLKBUF_X2 inst_11098 ( .A(net_9440), .Z(net_10946) );
AOI22_X2 inst_8226 ( .B1(net_8722), .A1(net_8500), .B2(net_4350), .A2(net_4349), .ZN(net_3811) );
CLKBUF_X2 inst_10706 ( .A(net_10553), .Z(net_10554) );
INV_X2 inst_6228 ( .ZN(net_5482), .A(net_5314) );
CLKBUF_X2 inst_15877 ( .A(net_15073), .Z(net_15725) );
INV_X4 inst_5236 ( .ZN(net_4889), .A(net_2580) );
CLKBUF_X2 inst_16602 ( .A(net_16449), .Z(net_16450) );
INV_X4 inst_5357 ( .ZN(net_1467), .A(net_1148) );
CLKBUF_X2 inst_12992 ( .A(net_12839), .Z(net_12840) );
CLKBUF_X2 inst_14204 ( .A(net_9301), .Z(net_14052) );
CLKBUF_X2 inst_16001 ( .A(net_13893), .Z(net_15849) );
CLKBUF_X2 inst_14104 ( .A(net_13951), .Z(net_13952) );
CLKBUF_X2 inst_9467 ( .A(net_9314), .Z(net_9315) );
CLKBUF_X2 inst_18277 ( .A(net_18124), .Z(net_18125) );
CLKBUF_X2 inst_17403 ( .A(net_10161), .Z(net_17251) );
CLKBUF_X2 inst_12231 ( .A(net_9945), .Z(net_12079) );
SDFFR_X1 inst_2682 ( .SI(net_7528), .SE(net_5043), .CK(net_11948), .RN(x6501), .Q(x4204), .D(x4204) );
AOI22_X2 inst_8517 ( .B1(net_6750), .A1(net_6717), .B2(net_6202), .A2(net_3520), .ZN(net_3423) );
CLKBUF_X2 inst_12434 ( .A(net_11688), .Z(net_12282) );
NAND2_X2 inst_4699 ( .A1(net_2931), .ZN(net_1882), .A2(net_1712) );
CLKBUF_X2 inst_10023 ( .A(net_9509), .Z(net_9871) );
NAND2_X2 inst_4749 ( .ZN(net_2704), .A1(net_1779), .A2(net_1586) );
SDFF_X2 inst_964 ( .SI(net_7322), .Q(net_6729), .D(net_6729), .SE(net_3124), .CK(net_9169) );
CLKBUF_X2 inst_16772 ( .A(net_16619), .Z(net_16620) );
NOR2_X2 inst_3372 ( .ZN(net_5553), .A1(net_5340), .A2(net_5339) );
AOI22_X2 inst_7940 ( .A1(net_7953), .B1(net_7783), .A2(net_6092), .B2(net_6091), .ZN(net_4185) );
CLKBUF_X2 inst_10165 ( .A(net_9271), .Z(net_10013) );
SDFFR_X2 inst_2313 ( .SE(net_2260), .Q(net_357), .D(net_357), .CK(net_11518), .RN(x6501), .SI(x2041) );
INV_X2 inst_6422 ( .ZN(net_756), .A(net_755) );
CLKBUF_X2 inst_10649 ( .A(net_10496), .Z(net_10497) );
CLKBUF_X2 inst_14778 ( .A(net_14625), .Z(net_14626) );
CLKBUF_X2 inst_12660 ( .A(net_11499), .Z(net_12508) );
CLKBUF_X2 inst_12629 ( .A(net_12476), .Z(net_12477) );
CLKBUF_X2 inst_14030 ( .A(net_13877), .Z(net_13878) );
CLKBUF_X2 inst_12965 ( .A(net_10943), .Z(net_12813) );
INV_X4 inst_6114 ( .ZN(net_1914), .A(net_263) );
CLKBUF_X2 inst_15359 ( .A(net_13486), .Z(net_15207) );
INV_X2 inst_6193 ( .A(net_6788), .ZN(net_5733) );
OAI21_X2 inst_3001 ( .B2(net_5902), .ZN(net_5892), .A(net_5816), .B1(net_770) );
CLKBUF_X2 inst_18032 ( .A(net_17879), .Z(net_17880) );
CLKBUF_X2 inst_14111 ( .A(net_11294), .Z(net_13959) );
CLKBUF_X2 inst_13741 ( .A(net_13588), .Z(net_13589) );
OR2_X4 inst_2818 ( .ZN(net_4396), .A2(net_4393), .A1(net_4369) );
OAI211_X2 inst_3198 ( .C1(net_8953), .ZN(net_2572), .C2(net_2466), .B(net_2394), .A(net_1310) );
CLKBUF_X2 inst_15893 ( .A(net_15740), .Z(net_15741) );
AOI22_X2 inst_7979 ( .B1(net_8196), .A1(net_7686), .B2(net_6099), .A2(net_4399), .ZN(net_4151) );
OAI33_X1 inst_2904 ( .A2(net_6416), .ZN(net_3150), .B3(net_3149), .A3(net_3149), .A1(net_2992), .B2(net_2991), .B1(net_1128) );
CLKBUF_X2 inst_10075 ( .A(net_9922), .Z(net_9923) );
CLKBUF_X2 inst_19092 ( .A(net_18595), .Z(net_18940) );
SDFFR_X2 inst_2383 ( .SI(net_7409), .SE(net_2260), .Q(net_346), .D(net_346), .CK(net_9361), .RN(x6501) );
SDFF_X2 inst_1701 ( .SI(net_7756), .Q(net_7756), .D(net_2590), .SE(net_2560), .CK(net_15967) );
CLKBUF_X2 inst_16933 ( .A(net_9945), .Z(net_16781) );
CLKBUF_X2 inst_12853 ( .A(net_12700), .Z(net_12701) );
CLKBUF_X2 inst_13853 ( .A(net_13700), .Z(net_13701) );
CLKBUF_X2 inst_10401 ( .A(net_10248), .Z(net_10249) );
CLKBUF_X2 inst_13577 ( .A(net_13424), .Z(net_13425) );
MUX2_X2 inst_4987 ( .A(net_9015), .Z(net_3961), .B(net_1457), .S(net_622) );
CLKBUF_X2 inst_9667 ( .A(net_9514), .Z(net_9515) );
CLKBUF_X2 inst_12262 ( .A(net_12109), .Z(net_12110) );
CLKBUF_X2 inst_9838 ( .A(net_9685), .Z(net_9686) );
CLKBUF_X2 inst_9627 ( .A(net_9118), .Z(net_9475) );
AND2_X2 inst_9163 ( .ZN(net_2828), .A1(net_2752), .A2(net_2751) );
CLKBUF_X2 inst_13405 ( .A(net_13252), .Z(net_13253) );
AOI222_X2 inst_8593 ( .ZN(net_3602), .A2(net_3599), .B2(net_3598), .C2(net_3597), .C1(net_3595), .B1(net_2089), .A1(net_1229) );
CLKBUF_X2 inst_14899 ( .A(net_14746), .Z(net_14747) );
DFFR_X2 inst_7228 ( .Q(net_6820), .D(net_2284), .CK(net_15190), .RN(x6501) );
CLKBUF_X2 inst_12503 ( .A(net_11322), .Z(net_12351) );
CLKBUF_X2 inst_9671 ( .A(net_9518), .Z(net_9519) );
SDFF_X2 inst_1135 ( .D(net_7310), .SI(net_6585), .Q(net_6585), .SE(net_3070), .CK(net_11864) );
AOI22_X2 inst_8333 ( .B1(net_8699), .A1(net_8662), .ZN(net_6222), .B2(net_6109), .A2(net_3857) );
CLKBUF_X2 inst_11871 ( .A(net_11718), .Z(net_11719) );
CLKBUF_X2 inst_14419 ( .A(net_13650), .Z(net_14267) );
OAI21_X2 inst_3127 ( .ZN(net_2215), .A(net_1966), .B2(net_1838), .B1(net_1648) );
CLKBUF_X2 inst_10945 ( .A(net_9981), .Z(net_10793) );
AOI221_X2 inst_8822 ( .B1(net_8984), .C2(net_5538), .B2(net_5456), .A(net_4898), .ZN(net_4582), .C1(net_413) );
CLKBUF_X2 inst_17595 ( .A(net_17442), .Z(net_17443) );
NOR4_X2 inst_3243 ( .ZN(net_1587), .A4(net_1038), .A1(net_1012), .A2(net_974), .A3(net_840) );
CLKBUF_X2 inst_14039 ( .A(net_13886), .Z(net_13887) );
AOI222_X1 inst_8605 ( .B2(net_6776), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5819), .A1(net_3116), .C1(x2746) );
CLKBUF_X2 inst_10564 ( .A(net_9850), .Z(net_10412) );
SDFF_X2 inst_1266 ( .Q(net_8084), .D(net_8084), .SI(net_2708), .SE(net_2707), .CK(net_15559) );
AOI21_X2 inst_8904 ( .ZN(net_5861), .A(net_5746), .B2(net_5661), .B1(net_4787) );
INV_X4 inst_5102 ( .ZN(net_5685), .A(net_5605) );
NAND2_X2 inst_4872 ( .A1(net_2549), .ZN(net_1072), .A2(net_807) );
CLKBUF_X2 inst_15781 ( .A(net_15628), .Z(net_15629) );
DFFR_X2 inst_7216 ( .QN(net_7361), .D(net_2380), .CK(net_11828), .RN(x6501) );
INV_X2 inst_6287 ( .ZN(net_4212), .A(net_3920) );
NAND2_X2 inst_4317 ( .A1(net_7138), .A2(net_5166), .ZN(net_5140) );
CLKBUF_X2 inst_13310 ( .A(net_12414), .Z(net_13158) );
DFFR_X2 inst_7090 ( .QN(net_8290), .D(net_3554), .CK(net_12062), .RN(x6501) );
CLKBUF_X2 inst_11379 ( .A(net_9211), .Z(net_11227) );
SDFF_X2 inst_1838 ( .D(net_7279), .SI(net_6896), .Q(net_6896), .SE(net_6284), .CK(net_14623) );
CLKBUF_X2 inst_9414 ( .A(net_9261), .Z(net_9262) );
SDFF_X2 inst_1454 ( .SI(net_7272), .Q(net_7089), .D(net_7089), .SE(net_6278), .CK(net_16846) );
CLKBUF_X2 inst_9438 ( .A(net_9198), .Z(net_9286) );
OAI21_X2 inst_3147 ( .A(net_2762), .B2(net_2250), .ZN(net_2005), .B1(net_1486) );
SDFF_X2 inst_1945 ( .SI(net_8049), .Q(net_8049), .D(net_2659), .SE(net_2508), .CK(net_18514) );
CLKBUF_X2 inst_16643 ( .A(net_16490), .Z(net_16491) );
INV_X4 inst_5564 ( .ZN(net_1521), .A(net_669) );
SDFFR_X1 inst_2657 ( .D(net_6779), .SE(net_4506), .CK(net_9185), .RN(x6501), .SI(x1500), .Q(x1500) );
INV_X4 inst_5722 ( .A(net_7241), .ZN(net_1945) );
CLKBUF_X2 inst_14581 ( .A(net_10361), .Z(net_14429) );
CLKBUF_X2 inst_13239 ( .A(net_13086), .Z(net_13087) );
CLKBUF_X2 inst_13043 ( .A(net_9714), .Z(net_12891) );
CLKBUF_X2 inst_12930 ( .A(net_12777), .Z(net_12778) );
SDFF_X2 inst_376 ( .SI(net_8376), .Q(net_8376), .SE(net_3969), .D(net_3965), .CK(net_10778) );
CLKBUF_X2 inst_10816 ( .A(net_10663), .Z(net_10664) );
CLKBUF_X2 inst_15356 ( .A(net_15203), .Z(net_15204) );
NOR3_X2 inst_3268 ( .A1(net_7308), .A2(net_6106), .ZN(net_2657), .A3(net_2449) );
CLKBUF_X2 inst_14066 ( .A(net_13913), .Z(net_13914) );
CLKBUF_X2 inst_17877 ( .A(net_17724), .Z(net_17725) );
CLKBUF_X2 inst_11676 ( .A(net_11523), .Z(net_11524) );
CLKBUF_X2 inst_14840 ( .A(net_9825), .Z(net_14688) );
CLKBUF_X2 inst_12167 ( .A(net_9601), .Z(net_12015) );
AOI22_X2 inst_7856 ( .A2(net_5595), .B2(net_5538), .ZN(net_4651), .B1(net_402), .A1(net_308) );
CLKBUF_X2 inst_10991 ( .A(net_10838), .Z(net_10839) );
AOI21_X2 inst_8897 ( .ZN(net_5786), .A(net_5785), .B2(net_5784), .B1(net_2668) );
INV_X2 inst_6299 ( .ZN(net_4042), .A(net_3908) );
CLKBUF_X2 inst_18250 ( .A(net_11641), .Z(net_18098) );
CLKBUF_X2 inst_12627 ( .A(net_12474), .Z(net_12475) );
CLKBUF_X2 inst_13251 ( .A(net_12311), .Z(net_13099) );
CLKBUF_X2 inst_10852 ( .A(net_9569), .Z(net_10700) );
CLKBUF_X2 inst_9951 ( .A(net_9798), .Z(net_9799) );
NAND3_X4 inst_3880 ( .A3(net_6085), .ZN(net_1562), .A1(net_1561), .A2(net_676) );
OAI21_X2 inst_3100 ( .ZN(net_2763), .A(net_2762), .B2(net_2506), .B1(net_2250) );
AOI22_X2 inst_8359 ( .B1(net_8702), .A1(net_8665), .B2(net_6109), .A2(net_3857), .ZN(net_3689) );
NAND2_X4 inst_4052 ( .ZN(net_6164), .A2(net_1662), .A1(net_1430) );
AOI22_X2 inst_8552 ( .B2(net_4889), .A1(net_4803), .ZN(net_3112), .B1(net_3111), .A2(net_2977) );
NAND2_X2 inst_4251 ( .A1(net_6908), .A2(net_5247), .ZN(net_5209) );
NAND2_X2 inst_4487 ( .A2(net_5609), .ZN(net_4485), .A1(net_362) );
SDFF_X2 inst_1596 ( .Q(net_8131), .D(net_8131), .SI(net_2722), .SE(net_2541), .CK(net_17696) );
NAND2_X2 inst_4364 ( .A1(net_7071), .A2(net_5162), .ZN(net_5093) );
CLKBUF_X2 inst_15313 ( .A(net_15160), .Z(net_15161) );
CLKBUF_X2 inst_15788 ( .A(net_15635), .Z(net_15636) );
INV_X2 inst_6400 ( .ZN(net_1154), .A(net_1153) );
DFFR_X2 inst_7078 ( .QN(net_7647), .D(net_3898), .CK(net_12695), .RN(x6501) );
CLKBUF_X2 inst_17145 ( .A(net_12092), .Z(net_16993) );
CLKBUF_X2 inst_10174 ( .A(net_10021), .Z(net_10022) );
SDFFR_X2 inst_2265 ( .D(net_7382), .SE(net_2797), .SI(net_191), .Q(net_191), .CK(net_14972), .RN(x6501) );
CLKBUF_X2 inst_13494 ( .A(net_13341), .Z(net_13342) );
SDFF_X2 inst_1555 ( .Q(net_7983), .D(net_7983), .SI(net_2658), .SE(net_2542), .CK(net_18054) );
SDFF_X2 inst_1293 ( .Q(net_8079), .D(net_8079), .SE(net_2707), .SI(net_2585), .CK(net_15777) );
DFFR_X2 inst_7132 ( .QN(net_5979), .D(net_3020), .CK(net_11222), .RN(x6501) );
NAND4_X2 inst_3805 ( .ZN(net_3621), .A1(net_3467), .A2(net_3466), .A3(net_3465), .A4(net_3464) );
XNOR2_X2 inst_280 ( .B(net_7374), .ZN(net_1025), .A(net_513) );
CLKBUF_X2 inst_11249 ( .A(net_9865), .Z(net_11097) );
OAI21_X2 inst_3157 ( .B2(net_2048), .ZN(net_1973), .A(net_1972), .B1(net_1691) );
CLKBUF_X2 inst_9888 ( .A(net_9147), .Z(net_9736) );
CLKBUF_X2 inst_11657 ( .A(net_11504), .Z(net_11505) );
CLKBUF_X2 inst_13648 ( .A(net_12556), .Z(net_13496) );
NAND2_X2 inst_4676 ( .ZN(net_2649), .A2(net_1924), .A1(net_1098) );
CLKBUF_X2 inst_17340 ( .A(net_17187), .Z(net_17188) );
CLKBUF_X2 inst_16958 ( .A(net_13164), .Z(net_16806) );
CLKBUF_X2 inst_14071 ( .A(net_13918), .Z(net_13919) );
CLKBUF_X2 inst_19129 ( .A(net_18976), .Z(net_18977) );
CLKBUF_X2 inst_16729 ( .A(net_16576), .Z(net_16577) );
AOI22_X2 inst_8110 ( .B1(net_8043), .A1(net_8009), .B2(net_6102), .A2(net_6097), .ZN(net_4037) );
CLKBUF_X2 inst_11556 ( .A(net_11403), .Z(net_11404) );
CLKBUF_X2 inst_14789 ( .A(net_14636), .Z(net_14637) );
CLKBUF_X2 inst_10344 ( .A(net_10043), .Z(net_10192) );
INV_X2 inst_6586 ( .A(net_6094), .ZN(net_6093) );
CLKBUF_X2 inst_15332 ( .A(net_12995), .Z(net_15180) );
CLKBUF_X2 inst_11188 ( .A(net_9416), .Z(net_11036) );
CLKBUF_X2 inst_17284 ( .A(net_17131), .Z(net_17132) );
NAND2_X2 inst_4393 ( .A1(net_7084), .A2(net_5164), .ZN(net_5064) );
AOI22_X2 inst_8299 ( .B1(net_8880), .A1(net_8325), .B2(net_6252), .A2(net_4345), .ZN(net_3744) );
CLKBUF_X2 inst_12743 ( .A(net_12590), .Z(net_12591) );
CLKBUF_X2 inst_17677 ( .A(net_17524), .Z(net_17525) );
CLKBUF_X2 inst_14780 ( .A(net_12133), .Z(net_14628) );
CLKBUF_X2 inst_18348 ( .A(net_16120), .Z(net_18196) );
SDFF_X2 inst_1359 ( .SI(net_7750), .Q(net_7750), .D(net_2574), .SE(net_2560), .CK(net_16069) );
CLKBUF_X2 inst_10345 ( .A(net_10192), .Z(net_10193) );
DFFR_X1 inst_7499 ( .Q(net_7300), .D(net_2256), .CK(net_15938), .RN(x6501) );
CLKBUF_X2 inst_14522 ( .A(net_14369), .Z(net_14370) );
CLKBUF_X2 inst_17209 ( .A(net_17056), .Z(net_17057) );
CLKBUF_X2 inst_11328 ( .A(net_9733), .Z(net_11176) );
NAND4_X2 inst_3797 ( .ZN(net_3629), .A1(net_3495), .A2(net_3494), .A3(net_3493), .A4(net_3492) );
XOR2_X1 inst_100 ( .A(net_6459), .B(net_3032), .Z(net_1214) );
NAND2_X2 inst_4352 ( .A1(net_7068), .A2(net_5162), .ZN(net_5105) );
XNOR2_X2 inst_279 ( .A(net_6365), .ZN(net_1027), .B(net_1026) );
CLKBUF_X2 inst_18468 ( .A(net_18315), .Z(net_18316) );
NOR2_X2 inst_3387 ( .A2(net_8220), .A1(net_4954), .ZN(net_4683) );
CLKBUF_X2 inst_11683 ( .A(net_11530), .Z(net_11531) );
CLKBUF_X2 inst_11014 ( .A(net_10861), .Z(net_10862) );
AOI22_X2 inst_8271 ( .B1(net_8876), .A1(net_8321), .B2(net_6252), .A2(net_4345), .ZN(net_3768) );
XOR2_X1 inst_81 ( .B(net_3272), .Z(net_3109), .A(net_2976) );
INV_X4 inst_5806 ( .A(net_8254), .ZN(net_542) );
CLKBUF_X2 inst_13424 ( .A(net_13271), .Z(net_13272) );
CLKBUF_X2 inst_9761 ( .A(net_9608), .Z(net_9609) );
DFFR_X2 inst_7087 ( .QN(net_7663), .D(net_3894), .CK(net_12672), .RN(x6501) );
CLKBUF_X2 inst_9471 ( .A(net_9318), .Z(net_9319) );
CLKBUF_X2 inst_14411 ( .A(net_14258), .Z(net_14259) );
CLKBUF_X2 inst_12040 ( .A(net_11887), .Z(net_11888) );
OAI221_X2 inst_2954 ( .ZN(net_4925), .C1(net_4924), .C2(net_4514), .B2(net_4475), .B1(net_2892), .A(net_2080) );
CLKBUF_X2 inst_9711 ( .A(net_9558), .Z(net_9559) );
CLKBUF_X2 inst_12045 ( .A(net_11892), .Z(net_11893) );
CLKBUF_X2 inst_11844 ( .A(net_11691), .Z(net_11692) );
SDFFR_X2 inst_2197 ( .SE(net_2517), .Q(net_304), .D(net_304), .SI(net_258), .CK(net_16425), .RN(x6501) );
AOI22_X2 inst_7995 ( .B1(net_8097), .A1(net_7757), .B2(net_6108), .A2(net_6096), .ZN(net_4138) );
CLKBUF_X2 inst_13064 ( .A(net_12911), .Z(net_12912) );
SDFFR_X2 inst_2582 ( .SI(net_7261), .Q(net_7261), .D(net_1461), .SE(net_1379), .CK(net_15027), .RN(x6501) );
XNOR2_X2 inst_142 ( .ZN(net_2303), .B(net_2232), .A(net_2231) );
XOR2_X1 inst_78 ( .B(net_3544), .Z(net_3235), .A(net_3105) );
CLKBUF_X2 inst_13182 ( .A(net_13029), .Z(net_13030) );
AOI22_X2 inst_7896 ( .B1(net_8978), .A2(net_5538), .B2(net_5456), .ZN(net_4533), .A1(net_407) );
OR3_X2 inst_2813 ( .ZN(net_1565), .A3(net_1304), .A1(net_552), .A2(x13921) );
XNOR2_X2 inst_177 ( .ZN(net_1734), .A(net_1463), .B(net_1238) );
SDFF_X2 inst_783 ( .SI(net_8353), .Q(net_8353), .D(net_3974), .SE(net_3880), .CK(net_10821) );
AOI22_X2 inst_7910 ( .A2(net_4553), .ZN(net_4514), .A1(net_4513), .B2(net_2066), .B1(net_1813) );
AOI22_X2 inst_8450 ( .B1(net_6735), .A1(net_6702), .B2(net_6202), .A2(net_3520), .ZN(net_3490) );
INV_X4 inst_5696 ( .ZN(net_628), .A(net_341) );
SDFF_X2 inst_2014 ( .SI(net_7927), .Q(net_7927), .D(net_2722), .SE(net_2461), .CK(net_17651) );
CLKBUF_X2 inst_14610 ( .A(net_14457), .Z(net_14458) );
INV_X4 inst_6122 ( .A(net_7218), .ZN(net_2981) );
CLKBUF_X2 inst_10144 ( .A(net_9991), .Z(net_9992) );
CLKBUF_X2 inst_12821 ( .A(net_12668), .Z(net_12669) );
CLKBUF_X2 inst_9999 ( .A(net_9822), .Z(net_9847) );
OR2_X4 inst_2822 ( .A1(net_4391), .ZN(net_4382), .A2(net_4370) );
SDFFR_X2 inst_2467 ( .SE(net_2260), .Q(net_365), .D(net_365), .CK(net_11447), .RN(x6501), .SI(x1804) );
INV_X2 inst_6176 ( .ZN(net_5914), .A(net_5867) );
CLKBUF_X2 inst_10335 ( .A(net_9411), .Z(net_10183) );
AOI222_X1 inst_8656 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3910), .B1(net_1764), .C1(net_1763), .A1(x13870) );
SDFF_X2 inst_2031 ( .SI(net_7780), .Q(net_7780), .D(net_2702), .SE(net_2459), .CK(net_18836) );
CLKBUF_X2 inst_18471 ( .A(net_18318), .Z(net_18319) );
NAND2_X2 inst_4386 ( .A1(net_7159), .A2(net_5166), .ZN(net_5071) );
CLKBUF_X2 inst_15367 ( .A(net_15060), .Z(net_15215) );
CLKBUF_X2 inst_14797 ( .A(net_14644), .Z(net_14645) );
CLKBUF_X2 inst_11282 ( .A(net_11129), .Z(net_11130) );
CLKBUF_X2 inst_16839 ( .A(net_16686), .Z(net_16687) );
CLKBUF_X2 inst_11527 ( .A(net_11374), .Z(net_11375) );
AOI22_X2 inst_8525 ( .B1(net_6722), .A1(net_6689), .B2(net_6202), .A2(net_3520), .ZN(net_3415) );
CLKBUF_X2 inst_17937 ( .A(net_17784), .Z(net_17785) );
XNOR2_X2 inst_338 ( .B(net_7393), .A(net_6375), .ZN(net_784) );
CLKBUF_X2 inst_16077 ( .A(net_15924), .Z(net_15925) );
INV_X4 inst_5577 ( .A(net_6371), .ZN(net_778) );
NAND3_X2 inst_4005 ( .ZN(net_1366), .A1(net_1266), .A3(net_1092), .A2(net_1084) );
INV_X4 inst_5424 ( .ZN(net_1126), .A(net_854) );
NAND2_X2 inst_4323 ( .A1(net_7121), .A2(net_5166), .ZN(net_5134) );
CLKBUF_X2 inst_17235 ( .A(net_17082), .Z(net_17083) );
CLKBUF_X2 inst_15212 ( .A(net_15059), .Z(net_15060) );
INV_X2 inst_6468 ( .ZN(net_2352), .A(net_157) );
CLKBUF_X2 inst_17397 ( .A(net_17244), .Z(net_17245) );
SDFFR_X2 inst_2474 ( .D(net_4697), .SE(net_2685), .SI(net_406), .Q(net_406), .CK(net_16649), .RN(x6501) );
SDFF_X2 inst_579 ( .Q(net_8845), .D(net_8845), .SE(net_3964), .SI(net_3940), .CK(net_10263) );
INV_X4 inst_5247 ( .ZN(net_2163), .A(net_1874) );
DFFR_X1 inst_7462 ( .D(net_4680), .CK(net_9588), .RN(x6501), .Q(x1130) );
SDFF_X2 inst_698 ( .Q(net_8440), .D(net_8440), .SI(net_3950), .SE(net_3934), .CK(net_12531) );
CLKBUF_X2 inst_14378 ( .A(net_14225), .Z(net_14226) );
NAND3_X2 inst_3964 ( .ZN(net_2510), .A1(net_2423), .A3(net_2402), .A2(net_2401) );
NAND3_X2 inst_3944 ( .ZN(net_4470), .A2(net_4469), .A3(net_4468), .A1(net_4275) );
NOR2_X2 inst_3394 ( .ZN(net_4491), .A2(net_4367), .A1(net_3929) );
CLKBUF_X2 inst_17280 ( .A(net_17127), .Z(net_17128) );
CLKBUF_X2 inst_17716 ( .A(net_17563), .Z(net_17564) );
INV_X4 inst_5978 ( .A(net_7229), .ZN(net_1806) );
OR2_X4 inst_2863 ( .ZN(net_6284), .A2(net_2199), .A1(net_1921) );
AOI22_X2 inst_8401 ( .B1(net_8822), .A1(net_8341), .A2(net_6265), .B2(net_6253), .ZN(net_3651) );
CLKBUF_X2 inst_12882 ( .A(net_12729), .Z(net_12730) );
CLKBUF_X2 inst_15565 ( .A(net_15403), .Z(net_15413) );
NAND3_X2 inst_3897 ( .ZN(net_5641), .A1(net_5570), .A3(net_5504), .A2(net_5406) );
INV_X4 inst_5534 ( .ZN(net_821), .A(net_655) );
CLKBUF_X2 inst_15897 ( .A(net_15744), .Z(net_15745) );
CLKBUF_X2 inst_11458 ( .A(net_11305), .Z(net_11306) );
CLKBUF_X2 inst_11693 ( .A(net_11540), .Z(net_11541) );
NAND4_X2 inst_3754 ( .A3(net_6073), .A1(net_6072), .ZN(net_4267), .A2(net_3871), .A4(net_3870) );
INV_X4 inst_6160 ( .A(net_6346), .ZN(net_6206) );
CLKBUF_X2 inst_15419 ( .A(net_15266), .Z(net_15267) );
CLKBUF_X2 inst_10229 ( .A(net_10076), .Z(net_10077) );
SDFF_X2 inst_837 ( .SI(net_8647), .Q(net_8647), .D(net_3967), .SE(net_3885), .CK(net_12416) );
INV_X4 inst_5716 ( .A(net_8296), .ZN(net_3550) );
CLKBUF_X2 inst_14425 ( .A(net_14272), .Z(net_14273) );
AOI21_X2 inst_8956 ( .A(net_5746), .ZN(net_5600), .B1(net_5259), .B2(net_5254) );
INV_X2 inst_6509 ( .A(net_7576), .ZN(net_3141) );
INV_X4 inst_5457 ( .ZN(net_2764), .A(net_1499) );
DFFR_X2 inst_7025 ( .QN(net_6305), .D(net_5694), .CK(net_16931), .RN(x6501) );
CLKBUF_X2 inst_14997 ( .A(net_12617), .Z(net_14845) );
AOI221_X2 inst_8785 ( .C2(net_6129), .B2(net_5609), .ZN(net_5038), .A(net_5022), .C1(net_1385), .B1(net_374) );
AOI22_X2 inst_7798 ( .A2(net_6130), .B2(net_4965), .ZN(net_4791), .A1(net_1421), .B1(net_387) );
CLKBUF_X2 inst_10497 ( .A(net_10344), .Z(net_10345) );
XOR2_X2 inst_65 ( .B(net_1033), .Z(net_923), .A(net_922) );
CLKBUF_X2 inst_12443 ( .A(net_12290), .Z(net_12291) );
CLKBUF_X2 inst_9563 ( .A(net_9375), .Z(net_9411) );
NOR2_X2 inst_3592 ( .A1(net_7353), .ZN(net_1269), .A2(net_1268) );
DFF_X1 inst_6822 ( .Q(net_8236), .D(net_4445), .CK(net_14454) );
INV_X4 inst_5121 ( .ZN(net_5463), .A(net_4471) );
NAND4_X2 inst_3732 ( .ZN(net_4298), .A1(net_4124), .A2(net_4123), .A3(net_4122), .A4(net_4121) );
CLKBUF_X2 inst_14931 ( .A(net_10531), .Z(net_14779) );
NAND2_X2 inst_4503 ( .A1(net_6273), .ZN(net_4376), .A2(net_1209) );
CLKBUF_X2 inst_9658 ( .A(net_9210), .Z(net_9506) );
NAND2_X2 inst_4907 ( .A2(net_7374), .ZN(net_610), .A1(net_163) );
OAI22_X2 inst_2926 ( .A2(net_2967), .B2(net_2943), .ZN(net_2891), .A1(net_2075), .B1(net_1323) );
CLKBUF_X2 inst_16392 ( .A(net_15684), .Z(net_16240) );
SDFF_X2 inst_1158 ( .SI(net_7313), .Q(net_6588), .D(net_6588), .SE(net_3069), .CK(net_11995) );
CLKBUF_X2 inst_18312 ( .A(net_18159), .Z(net_18160) );
AND2_X4 inst_9059 ( .A2(net_3325), .ZN(net_3319), .A1(net_3318) );
SDFF_X2 inst_1870 ( .D(net_7263), .SI(net_6960), .Q(net_6960), .SE(net_6283), .CK(net_14339) );
CLKBUF_X2 inst_13445 ( .A(net_13292), .Z(net_13293) );
DFFR_X2 inst_7038 ( .QN(net_7495), .D(net_4959), .CK(net_17254), .RN(x6501) );
INV_X4 inst_5270 ( .ZN(net_1871), .A(net_1782) );
CLKBUF_X2 inst_15853 ( .A(net_15700), .Z(net_15701) );
AOI22_X2 inst_8436 ( .B1(net_6533), .A1(net_6500), .A2(net_6137), .B2(net_6104), .ZN(net_3505) );
SDFFR_X2 inst_2445 ( .D(net_2916), .SE(net_2313), .SI(net_411), .Q(net_411), .CK(net_16660), .RN(x6501) );
CLKBUF_X2 inst_16205 ( .A(net_16052), .Z(net_16053) );
CLKBUF_X2 inst_14704 ( .A(net_14551), .Z(net_14552) );
OAI21_X2 inst_3039 ( .B2(net_8244), .B1(net_4928), .ZN(net_4831), .A(net_3200) );
INV_X4 inst_5477 ( .ZN(net_743), .A(net_742) );
CLKBUF_X2 inst_17277 ( .A(net_17124), .Z(net_17125) );
SDFF_X2 inst_461 ( .SI(net_8446), .Q(net_8446), .SE(net_3983), .D(net_3943), .CK(net_13361) );
INV_X4 inst_6092 ( .ZN(net_908), .A(net_186) );
AOI22_X2 inst_8291 ( .B1(net_8731), .A1(net_8509), .B2(net_4350), .A2(net_4349), .ZN(net_3751) );
INV_X2 inst_6387 ( .ZN(net_1303), .A(net_1302) );
SDFF_X2 inst_1973 ( .D(net_7268), .SI(net_6885), .Q(net_6885), .SE(net_6284), .CK(net_14312) );
OAI21_X2 inst_3051 ( .B2(net_8232), .B1(net_4850), .ZN(net_4760), .A(net_2613) );
AOI22_X2 inst_8326 ( .B1(net_8735), .A1(net_8513), .B2(net_4350), .A2(net_4349), .ZN(net_3720) );
SDFFR_X1 inst_2668 ( .D(net_6759), .SE(net_4506), .CK(net_11529), .RN(x6501), .SI(x2100), .Q(x2100) );
CLKBUF_X2 inst_14447 ( .A(net_14294), .Z(net_14295) );
CLKBUF_X2 inst_14238 ( .A(net_14085), .Z(net_14086) );
CLKBUF_X2 inst_17359 ( .A(net_17206), .Z(net_17207) );
INV_X4 inst_5742 ( .ZN(net_563), .A(x468) );
CLKBUF_X2 inst_18862 ( .A(net_18709), .Z(net_18710) );
INV_X4 inst_5775 ( .A(net_7421), .ZN(net_2462) );
NAND2_X2 inst_4808 ( .A2(net_2762), .ZN(net_1291), .A1(net_1290) );
NAND2_X2 inst_4657 ( .A1(net_2724), .A2(net_2334), .ZN(net_2271) );
SDFF_X2 inst_1669 ( .SI(net_7740), .Q(net_7740), .D(net_2705), .SE(net_2560), .CK(net_18537) );
DFFR_X1 inst_7456 ( .QN(net_8918), .D(net_4735), .CK(net_13964), .RN(x6501) );
CLKBUF_X2 inst_18973 ( .A(net_18820), .Z(net_18821) );
CLKBUF_X2 inst_17695 ( .A(net_17542), .Z(net_17543) );
CLKBUF_X2 inst_17690 ( .A(net_14723), .Z(net_17538) );
CLKBUF_X2 inst_12195 ( .A(net_9489), .Z(net_12043) );
CLKBUF_X2 inst_19082 ( .A(net_18929), .Z(net_18930) );
OAI21_X2 inst_3162 ( .ZN(net_2020), .A(net_1748), .B2(net_1439), .B1(net_1036) );
NAND3_X2 inst_3956 ( .ZN(net_3115), .A1(net_3114), .A2(net_2137), .A3(net_1489) );
SDFF_X2 inst_1801 ( .D(net_7276), .SI(net_6893), .Q(net_6893), .SE(net_6284), .CK(net_17372) );
CLKBUF_X2 inst_12777 ( .A(net_12624), .Z(net_12625) );
CLKBUF_X2 inst_9964 ( .A(net_9587), .Z(net_9812) );
SDFF_X2 inst_720 ( .SI(net_8516), .Q(net_8516), .D(net_3939), .SE(net_3884), .CK(net_10535) );
SDFF_X2 inst_958 ( .SI(net_7315), .Q(net_6689), .D(net_6689), .SE(net_3125), .CK(net_12137) );
CLKBUF_X2 inst_12412 ( .A(net_12259), .Z(net_12260) );
CLKBUF_X2 inst_10468 ( .A(net_10315), .Z(net_10316) );
CLKBUF_X2 inst_13465 ( .A(net_13235), .Z(net_13313) );
SDFF_X2 inst_368 ( .SI(net_8545), .Q(net_8545), .SE(net_3979), .D(net_3975), .CK(net_12563) );
SDFF_X2 inst_1697 ( .SI(net_7841), .Q(net_7841), .D(net_2585), .SE(net_2558), .CK(net_15749) );
CLKBUF_X2 inst_14909 ( .A(net_14756), .Z(net_14757) );
CLKBUF_X2 inst_14574 ( .A(net_14421), .Z(net_14422) );
DFFR_X2 inst_6995 ( .QN(net_6286), .D(net_5841), .CK(net_13883), .RN(x6501) );
CLKBUF_X2 inst_16269 ( .A(net_16116), .Z(net_16117) );
NAND4_X2 inst_3689 ( .ZN(net_4448), .A4(net_4348), .A1(net_3834), .A2(net_3833), .A3(net_3832) );
NOR2_X2 inst_3556 ( .A2(net_6169), .A1(net_6086), .ZN(net_1367) );
CLKBUF_X2 inst_17157 ( .A(net_16254), .Z(net_17005) );
CLKBUF_X2 inst_17670 ( .A(net_17517), .Z(net_17518) );
AOI221_X2 inst_8811 ( .C2(net_5609), .B2(net_5520), .A(net_4834), .ZN(net_4717), .C1(net_355), .B1(net_285) );
SDFF_X2 inst_1966 ( .D(net_7279), .SI(net_7016), .Q(net_7016), .SE(net_6277), .CK(net_14599) );
NAND3_X2 inst_3914 ( .ZN(net_5624), .A1(net_5553), .A3(net_5487), .A2(net_5338) );
NAND2_X2 inst_4716 ( .A1(net_2499), .ZN(net_1786), .A2(net_1783) );
DFF_X1 inst_6838 ( .Q(net_6428), .D(net_3609), .CK(net_17980) );
CLKBUF_X2 inst_18076 ( .A(net_17923), .Z(net_17924) );
SDFFR_X2 inst_2435 ( .D(net_3203), .SE(net_2313), .SI(net_423), .Q(net_423), .CK(net_14820), .RN(x6501) );
CLKBUF_X2 inst_17946 ( .A(net_17793), .Z(net_17794) );
CLKBUF_X2 inst_16673 ( .A(net_16520), .Z(net_16521) );
CLKBUF_X2 inst_14078 ( .A(net_13309), .Z(net_13926) );
CLKBUF_X2 inst_10101 ( .A(net_9948), .Z(net_9949) );
CLKBUF_X2 inst_18210 ( .A(net_18057), .Z(net_18058) );
SDFF_X2 inst_1678 ( .SI(net_7863), .Q(net_7863), .D(net_2749), .SE(net_2558), .CK(net_13759) );
CLKBUF_X2 inst_19169 ( .A(net_19016), .Z(net_19017) );
CLKBUF_X2 inst_11602 ( .A(net_11449), .Z(net_11450) );
CLKBUF_X2 inst_10839 ( .A(net_10686), .Z(net_10687) );
CLKBUF_X2 inst_15424 ( .A(net_13581), .Z(net_15272) );
SDFFR_X2 inst_2233 ( .Q(net_7467), .D(net_7467), .SE(net_2863), .CK(net_12161), .SI(x13457), .RN(x6501) );
CLKBUF_X2 inst_17033 ( .A(net_16880), .Z(net_16881) );
DFFR_X2 inst_7266 ( .QN(net_6380), .D(net_1995), .CK(net_18258), .RN(x6501) );
CLKBUF_X2 inst_14859 ( .A(net_14706), .Z(net_14707) );
CLKBUF_X2 inst_13939 ( .A(net_13786), .Z(net_13787) );
CLKBUF_X2 inst_13870 ( .A(net_13471), .Z(net_13718) );
SDFF_X2 inst_396 ( .SI(net_8307), .Q(net_8307), .SE(net_3978), .D(net_3960), .CK(net_13367) );
NOR2_X2 inst_3382 ( .ZN(net_5543), .A1(net_5297), .A2(net_5296) );
CLKBUF_X2 inst_15548 ( .A(net_10422), .Z(net_15396) );
NOR2_X2 inst_3377 ( .ZN(net_5548), .A1(net_5317), .A2(net_5316) );
INV_X4 inst_5128 ( .ZN(net_4468), .A(net_4406) );
CLKBUF_X2 inst_14665 ( .A(net_14512), .Z(net_14513) );
CLKBUF_X2 inst_14330 ( .A(net_10589), .Z(net_14178) );
CLKBUF_X2 inst_10371 ( .A(net_10218), .Z(net_10219) );
CLKBUF_X2 inst_11894 ( .A(net_11741), .Z(net_11742) );
CLKBUF_X2 inst_14992 ( .A(net_14839), .Z(net_14840) );
OR2_X4 inst_2845 ( .ZN(net_2248), .A2(net_2071), .A1(net_1663) );
AOI22_X2 inst_7760 ( .B1(net_6988), .A1(net_6948), .A2(net_5443), .B2(net_5442), .ZN(net_5366) );
OAI221_X2 inst_2977 ( .ZN(net_1460), .C2(net_1459), .A(net_794), .C1(net_679), .B2(net_678), .B1(net_634) );
SDFF_X2 inst_1092 ( .D(net_7317), .SI(net_6493), .Q(net_6493), .SE(net_3071), .CK(net_9850) );
CLKBUF_X2 inst_11181 ( .A(net_11028), .Z(net_11029) );
CLKBUF_X2 inst_9843 ( .A(net_9690), .Z(net_9691) );
DFFR_X1 inst_7492 ( .QN(net_6473), .D(net_3341), .CK(net_15136), .RN(x6501) );
CLKBUF_X2 inst_18962 ( .A(net_18809), .Z(net_18810) );
CLKBUF_X2 inst_11784 ( .A(net_11538), .Z(net_11632) );
CLKBUF_X2 inst_15729 ( .A(net_15576), .Z(net_15577) );
CLKBUF_X2 inst_19170 ( .A(net_18803), .Z(net_19018) );
CLKBUF_X2 inst_10011 ( .A(net_9858), .Z(net_9859) );
CLKBUF_X2 inst_14231 ( .A(net_14078), .Z(net_14079) );
CLKBUF_X2 inst_16637 ( .A(net_15319), .Z(net_16485) );
CLKBUF_X2 inst_16920 ( .A(net_16767), .Z(net_16768) );
CLKBUF_X2 inst_11356 ( .A(net_11130), .Z(net_11204) );
AOI22_X2 inst_7780 ( .A1(net_5268), .B2(net_5267), .ZN(net_4871), .A2(net_4635), .B1(net_178) );
NAND2_X2 inst_4592 ( .ZN(net_3927), .A1(net_2847), .A2(net_2846) );
CLKBUF_X2 inst_15696 ( .A(net_15543), .Z(net_15544) );
SDFF_X2 inst_451 ( .Q(net_8749), .D(net_8749), .SE(net_3982), .SI(net_3937), .CK(net_13058) );
INV_X4 inst_5478 ( .A(net_1568), .ZN(net_741) );
SDFFR_X2 inst_2166 ( .QN(net_7588), .D(net_3941), .SE(net_3144), .SI(net_3135), .CK(net_10395), .RN(x6501) );
CLKBUF_X2 inst_16145 ( .A(net_15992), .Z(net_15993) );
CLKBUF_X2 inst_14486 ( .A(net_11561), .Z(net_14334) );
CLKBUF_X2 inst_15377 ( .A(net_15224), .Z(net_15225) );
CLKBUF_X2 inst_9910 ( .A(net_9227), .Z(net_9758) );
DFFR_X1 inst_7471 ( .QN(net_7421), .D(net_4217), .CK(net_13386), .RN(x6501) );
DFFR_X2 inst_7221 ( .D(net_2372), .QN(net_215), .CK(net_17562), .RN(x6501) );
CLKBUF_X2 inst_18193 ( .A(net_18040), .Z(net_18041) );
INV_X4 inst_5295 ( .A(net_1814), .ZN(net_1600) );
NAND4_X2 inst_3657 ( .A4(net_6038), .A1(net_6037), .ZN(net_4608), .A2(net_4150), .A3(net_4149) );
DFFR_X2 inst_7319 ( .D(net_8288), .QN(net_8284), .CK(net_12224), .RN(x6501) );
DFFS_X2 inst_6896 ( .Q(net_7480), .D(net_2645), .CK(net_16151), .SN(x6501) );
CLKBUF_X2 inst_14529 ( .A(net_14376), .Z(net_14377) );
CLKBUF_X2 inst_17682 ( .A(net_17529), .Z(net_17530) );
SDFF_X2 inst_1998 ( .SI(net_7920), .Q(net_7920), .D(net_2574), .SE(net_2461), .CK(net_18347) );
CLKBUF_X2 inst_17382 ( .A(net_17229), .Z(net_17230) );
NOR3_X2 inst_3302 ( .A2(net_2843), .ZN(net_1800), .A1(net_1799), .A3(net_1499) );
CLKBUF_X2 inst_11157 ( .A(net_11004), .Z(net_11005) );
CLKBUF_X2 inst_16793 ( .A(net_16640), .Z(net_16641) );
OR2_X2 inst_2870 ( .ZN(net_5597), .A2(net_5454), .A1(net_3161) );
CLKBUF_X2 inst_14902 ( .A(net_14749), .Z(net_14750) );
SDFF_X2 inst_874 ( .Q(net_8585), .D(net_8585), .SI(net_3952), .SE(net_3878), .CK(net_12855) );
CLKBUF_X2 inst_17991 ( .A(net_15050), .Z(net_17839) );
SDFF_X2 inst_1681 ( .Q(net_8176), .D(net_8176), .SI(net_2704), .SE(net_2538), .CK(net_16989) );
CLKBUF_X2 inst_10222 ( .A(net_10069), .Z(net_10070) );
AND2_X2 inst_9173 ( .A1(net_2693), .ZN(net_2587), .A2(net_2483) );
SDFF_X2 inst_1652 ( .SI(net_7735), .Q(net_7735), .D(net_2716), .SE(net_2559), .CK(net_17064) );
CLKBUF_X2 inst_9391 ( .A(net_9238), .Z(net_9239) );
CLKBUF_X2 inst_15576 ( .A(net_15423), .Z(net_15424) );
SDFF_X2 inst_1622 ( .Q(net_8165), .D(net_8165), .SI(net_2722), .SE(net_2538), .CK(net_18782) );
CLKBUF_X2 inst_13965 ( .A(net_13812), .Z(net_13813) );
SDFF_X2 inst_1735 ( .SI(net_7292), .Q(net_7149), .D(net_7149), .SE(net_6279), .CK(net_14904) );
SDFF_X2 inst_2050 ( .SI(net_7919), .Q(net_7919), .D(net_2706), .SE(net_2461), .CK(net_15219) );
CLKBUF_X2 inst_9516 ( .A(net_9363), .Z(net_9364) );
INV_X4 inst_5458 ( .ZN(net_772), .A(net_771) );
NAND2_X2 inst_4555 ( .A1(net_6384), .A2(net_6184), .ZN(net_3255) );
CLKBUF_X2 inst_16366 ( .A(net_11876), .Z(net_16214) );
AOI222_X1 inst_8681 ( .B1(net_6754), .A1(net_6462), .C1(net_6459), .A2(net_3296), .B2(net_3295), .C2(net_3294), .ZN(net_3291) );
SDFF_X2 inst_1189 ( .D(net_7331), .SI(net_6573), .Q(net_6573), .SE(net_3070), .CK(net_11639) );
CLKBUF_X2 inst_15762 ( .A(net_15609), .Z(net_15610) );
SDFFR_X2 inst_2360 ( .SE(net_2260), .Q(net_309), .D(net_309), .CK(net_9309), .RN(x6501), .SI(x3561) );
CLKBUF_X2 inst_16847 ( .A(net_10908), .Z(net_16695) );
CLKBUF_X2 inst_11052 ( .A(net_10899), .Z(net_10900) );
CLKBUF_X2 inst_16460 ( .A(net_16307), .Z(net_16308) );
CLKBUF_X2 inst_16401 ( .A(net_16248), .Z(net_16249) );
XOR2_X2 inst_33 ( .A(net_2728), .B(net_2677), .Z(net_1192) );
SDFFR_X2 inst_2107 ( .SI(net_7407), .Q(net_7407), .SE(net_6198), .D(net_5733), .CK(net_9384), .RN(x6501) );
CLKBUF_X2 inst_12756 ( .A(net_12603), .Z(net_12604) );
XNOR2_X2 inst_232 ( .ZN(net_1297), .A(net_1296), .B(net_711) );
CLKBUF_X2 inst_16764 ( .A(net_9911), .Z(net_16612) );
INV_X2 inst_6253 ( .ZN(net_4846), .A(net_4737) );
DFFR_X1 inst_7575 ( .D(net_6482), .Q(net_6464), .CK(net_15122), .RN(x6501) );
NAND2_X2 inst_4628 ( .ZN(net_2892), .A2(net_2642), .A1(net_2528) );
CLKBUF_X2 inst_16452 ( .A(net_15590), .Z(net_16300) );
NAND4_X2 inst_3794 ( .ZN(net_3632), .A1(net_3512), .A2(net_3511), .A3(net_3510), .A4(net_3509) );
CLKBUF_X2 inst_9648 ( .A(net_9495), .Z(net_9496) );
CLKBUF_X2 inst_18904 ( .A(net_18751), .Z(net_18752) );
CLKBUF_X2 inst_18704 ( .A(net_11932), .Z(net_18552) );
CLKBUF_X2 inst_14463 ( .A(net_9719), .Z(net_14311) );
CLKBUF_X2 inst_16317 ( .A(net_12844), .Z(net_16165) );
CLKBUF_X2 inst_9608 ( .A(net_9455), .Z(net_9456) );
CLKBUF_X1 inst_7730 ( .A(x192486), .Z(x1024) );
CLKBUF_X2 inst_13945 ( .A(net_12995), .Z(net_13793) );
NAND4_X2 inst_3652 ( .A4(net_6000), .A1(net_5999), .ZN(net_4613), .A3(net_4180), .A2(net_4179) );
CLKBUF_X2 inst_12428 ( .A(net_12275), .Z(net_12276) );
CLKBUF_X2 inst_18185 ( .A(net_11933), .Z(net_18033) );
CLKBUF_X2 inst_14513 ( .A(net_13094), .Z(net_14361) );
INV_X8 inst_5043 ( .ZN(net_6107), .A(net_3572) );
CLKBUF_X2 inst_17635 ( .A(net_17482), .Z(net_17483) );
CLKBUF_X2 inst_18266 ( .A(net_12535), .Z(net_18114) );
CLKBUF_X2 inst_13751 ( .A(net_11631), .Z(net_13599) );
DFFS_X2 inst_6907 ( .QN(net_8268), .D(net_8264), .CK(net_18465), .SN(x6501) );
CLKBUF_X2 inst_9331 ( .A(net_9178), .Z(net_9179) );
SDFF_X2 inst_602 ( .SI(net_8396), .Q(net_8396), .SE(net_3969), .D(net_3954), .CK(net_10928) );
CLKBUF_X2 inst_18945 ( .A(net_18792), .Z(net_18793) );
XNOR2_X2 inst_135 ( .ZN(net_2746), .A(net_2554), .B(net_2551) );
CLKBUF_X2 inst_10091 ( .A(net_9938), .Z(net_9939) );
CLKBUF_X2 inst_11711 ( .A(net_11558), .Z(net_11559) );
CLKBUF_X2 inst_17705 ( .A(net_17108), .Z(net_17553) );
CLKBUF_X2 inst_10037 ( .A(net_9593), .Z(net_9885) );
CLKBUF_X2 inst_18241 ( .A(net_18088), .Z(net_18089) );
CLKBUF_X2 inst_9321 ( .A(net_9168), .Z(net_9169) );
OAI21_X2 inst_3117 ( .B1(net_6418), .ZN(net_2337), .A(net_2184), .B2(net_2183) );
CLKBUF_X2 inst_16763 ( .A(net_15360), .Z(net_16611) );
INV_X4 inst_6072 ( .A(net_7491), .ZN(net_754) );
NAND4_X2 inst_3770 ( .A3(net_6067), .A1(net_6066), .ZN(net_4251), .A2(net_3766), .A4(net_3765) );
AOI22_X2 inst_8157 ( .B1(net_8087), .A1(net_7747), .B2(net_6108), .A2(net_6096), .ZN(net_3995) );
CLKBUF_X2 inst_13863 ( .A(net_13710), .Z(net_13711) );
CLKBUF_X2 inst_16260 ( .A(net_12181), .Z(net_16108) );
SDFFR_X1 inst_2709 ( .SI(net_6813), .Q(net_6813), .D(net_6810), .SE(net_6270), .CK(net_11793), .RN(x6501) );
XNOR2_X2 inst_224 ( .ZN(net_1382), .B(net_1381), .A(net_616) );
CLKBUF_X2 inst_14756 ( .A(net_14603), .Z(net_14604) );
CLKBUF_X2 inst_14003 ( .A(net_13850), .Z(net_13851) );
CLKBUF_X2 inst_9661 ( .A(net_9508), .Z(net_9509) );
NAND4_X2 inst_3635 ( .ZN(net_5327), .A2(net_4968), .A4(net_4866), .A1(net_4805), .A3(net_4574) );
CLKBUF_X2 inst_16481 ( .A(net_12629), .Z(net_16329) );
INV_X4 inst_5399 ( .ZN(net_3535), .A(net_882) );
INV_X8 inst_5058 ( .ZN(net_6263), .A(net_3314) );
CLKBUF_X2 inst_14297 ( .A(net_9983), .Z(net_14145) );
SDFFR_X2 inst_2406 ( .D(net_7374), .SI(net_2692), .SE(net_2316), .QN(net_276), .CK(net_16415), .RN(x6501) );
AOI221_X2 inst_8796 ( .C2(net_6187), .B2(net_5609), .ZN(net_4899), .A(net_4898), .B1(net_373), .C1(net_197) );
CLKBUF_X2 inst_17994 ( .A(net_17841), .Z(net_17842) );
SDFF_X2 inst_801 ( .SI(net_8342), .Q(net_8342), .D(net_3937), .SE(net_3880), .CK(net_10704) );
CLKBUF_X2 inst_10617 ( .A(net_10351), .Z(net_10465) );
CLKBUF_X2 inst_16873 ( .A(net_12511), .Z(net_16721) );
SDFF_X2 inst_870 ( .Q(net_8580), .D(net_8580), .SI(net_3955), .SE(net_3878), .CK(net_10966) );
CLKBUF_X2 inst_12544 ( .A(net_9441), .Z(net_12392) );
CLKBUF_X2 inst_9660 ( .A(net_9251), .Z(net_9508) );
XOR2_X2 inst_11 ( .A(net_6800), .Z(net_1666), .B(net_1234) );
CLKBUF_X2 inst_15537 ( .A(net_15384), .Z(net_15385) );
CLKBUF_X2 inst_13468 ( .A(net_13315), .Z(net_13316) );
SDFFR_X2 inst_2276 ( .SI(net_7389), .SE(net_2814), .Q(net_248), .D(net_248), .CK(net_14709), .RN(x6501) );
AOI21_X2 inst_8892 ( .B2(net_5871), .ZN(net_5796), .A(net_5795), .B1(net_2667) );
SDFFR_X2 inst_2301 ( .D(net_3544), .SE(net_2748), .SI(net_414), .Q(net_414), .CK(net_17288), .RN(x6501) );
CLKBUF_X2 inst_18404 ( .A(net_18251), .Z(net_18252) );
AOI22_X2 inst_8202 ( .B1(net_8830), .A1(net_8349), .A2(net_6265), .B2(net_6253), .ZN(net_3834) );
SDFF_X2 inst_557 ( .Q(net_8671), .D(net_8671), .SI(net_3938), .SE(net_3935), .CK(net_12989) );
CLKBUF_X2 inst_13639 ( .A(net_13486), .Z(net_13487) );
CLKBUF_X2 inst_14300 ( .A(net_14147), .Z(net_14148) );
CLKBUF_X2 inst_11154 ( .A(net_9666), .Z(net_11002) );
NOR3_X2 inst_3279 ( .ZN(net_2795), .A1(net_2400), .A3(net_2396), .A2(net_1127) );
SDFF_X2 inst_823 ( .SI(net_8515), .Q(net_8515), .D(net_3976), .SE(net_3884), .CK(net_10323) );
SDFF_X2 inst_1461 ( .SI(net_7284), .Q(net_7141), .D(net_7141), .SE(net_6279), .CK(net_16220) );
AOI221_X2 inst_8809 ( .C2(net_5535), .B2(net_5260), .A(net_4898), .ZN(net_4719), .B1(net_3332), .C1(net_474) );
NAND4_X2 inst_3773 ( .ZN(net_4248), .A1(net_3748), .A2(net_3747), .A3(net_3746), .A4(net_3745) );
NAND2_X2 inst_4767 ( .ZN(net_4394), .A1(net_1802), .A2(net_1679) );
CLKBUF_X2 inst_10608 ( .A(net_10237), .Z(net_10456) );
CLKBUF_X2 inst_19014 ( .A(net_15802), .Z(net_18862) );
CLKBUF_X2 inst_13154 ( .A(net_12613), .Z(net_13002) );
INV_X4 inst_5620 ( .A(net_7378), .ZN(net_1023) );
CLKBUF_X2 inst_11409 ( .A(net_9061), .Z(net_11257) );
DFFR_X2 inst_7104 ( .QN(net_8259), .D(net_3207), .CK(net_18503), .RN(x6501) );
AOI22_X2 inst_7746 ( .B1(net_6975), .A1(net_6935), .A2(net_5443), .B2(net_5442), .ZN(net_5422) );
CLKBUF_X2 inst_9976 ( .A(net_9823), .Z(net_9824) );
AOI22_X2 inst_8342 ( .B1(net_8774), .A1(net_8404), .A2(net_3867), .B2(net_3866), .ZN(net_3705) );
CLKBUF_X2 inst_18121 ( .A(net_17968), .Z(net_17969) );
CLKBUF_X2 inst_14084 ( .A(net_13931), .Z(net_13932) );
CLKBUF_X2 inst_16544 ( .A(net_13299), .Z(net_16392) );
SDFF_X2 inst_1413 ( .Q(net_7076), .D(net_7076), .SE(net_6280), .SI(net_2544), .CK(net_15906) );
CLKBUF_X2 inst_13320 ( .A(net_13167), .Z(net_13168) );
NAND3_X2 inst_3993 ( .ZN(net_1748), .A1(net_1120), .A3(net_1030), .A2(net_991) );
DFFS_X1 inst_6926 ( .D(net_6145), .CK(net_16372), .SN(x6501), .Q(x831) );
CLKBUF_X2 inst_11140 ( .A(net_10987), .Z(net_10988) );
CLKBUF_X2 inst_17615 ( .A(net_17462), .Z(net_17463) );
CLKBUF_X2 inst_13272 ( .A(net_13119), .Z(net_13120) );
CLKBUF_X2 inst_16161 ( .A(net_12764), .Z(net_16009) );
SDFFR_X2 inst_2169 ( .QN(net_7565), .D(net_3938), .SE(net_3144), .SI(net_3133), .CK(net_10792), .RN(x6501) );
CLKBUF_X2 inst_11903 ( .A(net_9200), .Z(net_11751) );
CLKBUF_X2 inst_15258 ( .A(net_11710), .Z(net_15106) );
SDFF_X2 inst_1326 ( .SI(net_7685), .Q(net_7685), .SE(net_2714), .D(net_2576), .CK(net_16074) );
CLKBUF_X2 inst_18065 ( .A(net_11727), .Z(net_17913) );
AOI21_X2 inst_8960 ( .ZN(net_3882), .B2(net_3552), .B1(net_3550), .A(net_3362) );
CLKBUF_X2 inst_16473 ( .A(net_16320), .Z(net_16321) );
CLKBUF_X2 inst_14938 ( .A(net_14785), .Z(net_14786) );
AOI22_X2 inst_8191 ( .B1(net_8717), .A1(net_8495), .ZN(net_6075), .B2(net_4350), .A2(net_4349) );
CLKBUF_X2 inst_11920 ( .A(net_11767), .Z(net_11768) );
NAND2_X2 inst_4238 ( .A1(net_7022), .A2(net_5249), .ZN(net_5222) );
CLKBUF_X2 inst_9496 ( .A(net_9259), .Z(net_9344) );
INV_X4 inst_5275 ( .ZN(net_1687), .A(net_1686) );
CLKBUF_X2 inst_18029 ( .A(net_17876), .Z(net_17877) );
CLKBUF_X2 inst_18800 ( .A(net_12179), .Z(net_18648) );
CLKBUF_X2 inst_14791 ( .A(net_12287), .Z(net_14639) );
CLKBUF_X2 inst_14887 ( .A(net_10446), .Z(net_14735) );
CLKBUF_X2 inst_16374 ( .A(net_16221), .Z(net_16222) );
AND2_X2 inst_9197 ( .A1(net_7260), .ZN(net_6057), .A2(net_1377) );
INV_X4 inst_6127 ( .A(net_7376), .ZN(net_1118) );
CLKBUF_X2 inst_14867 ( .A(net_10199), .Z(net_14715) );
SDFFR_X2 inst_2154 ( .Q(net_8280), .D(net_3233), .SI(net_3029), .SE(net_2996), .CK(net_18440), .RN(x6501) );
CLKBUF_X2 inst_16487 ( .A(net_16334), .Z(net_16335) );
NAND2_X2 inst_4602 ( .ZN(net_2665), .A2(net_2664), .A1(net_2447) );
SDFFR_X2 inst_2602 ( .D(net_7371), .Q(net_7268), .SI(net_1855), .SE(net_1327), .CK(net_14682), .RN(x6501) );
XNOR2_X2 inst_109 ( .ZN(net_5019), .A(net_4705), .B(net_1538) );
SDFF_X2 inst_1182 ( .SI(net_7312), .Q(net_6587), .D(net_6587), .SE(net_3069), .CK(net_11990) );
DFFS_X2 inst_6875 ( .QN(net_7646), .D(net_3899), .CK(net_12664), .SN(x6501) );
NAND3_X2 inst_3983 ( .A2(net_7374), .A1(net_2315), .ZN(net_2292), .A3(net_1932) );
CLKBUF_X2 inst_15066 ( .A(net_14913), .Z(net_14914) );
CLKBUF_X2 inst_17311 ( .A(net_10942), .Z(net_17159) );
CLKBUF_X2 inst_12275 ( .A(net_9404), .Z(net_12123) );
CLKBUF_X2 inst_11019 ( .A(net_10646), .Z(net_10867) );
INV_X4 inst_5984 ( .A(net_6299), .ZN(net_2671) );
SDFF_X2 inst_1444 ( .SI(net_7290), .Q(net_7107), .D(net_7107), .SE(net_6278), .CK(net_18283) );
CLKBUF_X2 inst_11993 ( .A(net_11840), .Z(net_11841) );
INV_X4 inst_5490 ( .ZN(net_724), .A(net_723) );
CLKBUF_X2 inst_17226 ( .A(net_14133), .Z(net_17074) );
SDFF_X2 inst_1231 ( .Q(net_7823), .D(net_7823), .SE(net_2730), .SI(net_2719), .CK(net_15638) );
CLKBUF_X2 inst_15557 ( .A(net_15404), .Z(net_15405) );
SDFF_X2 inst_904 ( .SI(net_8722), .Q(net_8722), .SE(net_6195), .D(net_3958), .CK(net_12233) );
CLKBUF_X2 inst_12100 ( .A(net_11525), .Z(net_11948) );
CLKBUF_X2 inst_10628 ( .A(net_10475), .Z(net_10476) );
CLKBUF_X2 inst_13147 ( .A(net_12994), .Z(net_12995) );
SDFFR_X2 inst_2159 ( .QN(net_7576), .D(net_3973), .SE(net_3144), .SI(net_3141), .CK(net_10951), .RN(x6501) );
CLKBUF_X2 inst_18012 ( .A(net_17859), .Z(net_17860) );
DFFR_X2 inst_7051 ( .QN(net_7508), .D(net_4840), .CK(net_14837), .RN(x6501) );
INV_X2 inst_6266 ( .A(net_8248), .ZN(net_4631) );
NAND3_X2 inst_3923 ( .ZN(net_5615), .A1(net_5544), .A3(net_5478), .A2(net_5299) );
CLKBUF_X2 inst_16042 ( .A(net_15889), .Z(net_15890) );
NAND2_X2 inst_4831 ( .A1(net_6406), .A2(net_6405), .ZN(net_2909) );
SDFF_X2 inst_757 ( .Q(net_8798), .D(net_8798), .SI(net_3957), .SE(net_3879), .CK(net_10986) );
SDFF_X2 inst_1627 ( .Q(net_8171), .D(net_8171), .SI(net_2711), .SE(net_2538), .CK(net_14268) );
CLKBUF_X2 inst_18629 ( .A(net_9750), .Z(net_18477) );
CLKBUF_X2 inst_12670 ( .A(net_12517), .Z(net_12518) );
CLKBUF_X2 inst_17857 ( .A(net_17704), .Z(net_17705) );
CLKBUF_X2 inst_13557 ( .A(net_13404), .Z(net_13405) );
CLKBUF_X2 inst_12994 ( .A(net_9362), .Z(net_12842) );
NAND4_X2 inst_3817 ( .ZN(net_3609), .A1(net_3419), .A2(net_3418), .A3(net_3417), .A4(net_3416) );
CLKBUF_X2 inst_15201 ( .A(net_14966), .Z(net_15049) );
CLKBUF_X2 inst_15458 ( .A(net_15305), .Z(net_15306) );
INV_X4 inst_5065 ( .ZN(net_5915), .A(net_5868) );
SDFF_X2 inst_1256 ( .Q(net_8089), .D(net_8089), .SE(net_2707), .SI(net_2706), .CK(net_18898) );
CLKBUF_X2 inst_17204 ( .A(net_17051), .Z(net_17052) );
CLKBUF_X2 inst_15710 ( .A(net_15557), .Z(net_15558) );
CLKBUF_X2 inst_9549 ( .A(net_9396), .Z(net_9397) );
CLKBUF_X2 inst_15752 ( .A(net_15599), .Z(net_15600) );
SDFF_X2 inst_1903 ( .D(net_7301), .SI(net_7038), .Q(net_7038), .SE(net_6277), .CK(net_15871) );
CLKBUF_X2 inst_14254 ( .A(net_14101), .Z(net_14102) );
CLKBUF_X2 inst_9503 ( .A(net_9350), .Z(net_9351) );
CLKBUF_X2 inst_11230 ( .A(net_11077), .Z(net_11078) );
CLKBUF_X2 inst_13716 ( .A(net_13563), .Z(net_13564) );
SDFFR_X2 inst_2554 ( .QN(net_6370), .SE(net_2147), .SI(net_1946), .D(net_780), .CK(net_18133), .RN(x6501) );
CLKBUF_X2 inst_16993 ( .A(net_12253), .Z(net_16841) );
CLKBUF_X2 inst_9423 ( .A(net_9270), .Z(net_9271) );
CLKBUF_X2 inst_14422 ( .A(net_14269), .Z(net_14270) );
CLKBUF_X2 inst_15295 ( .A(net_15142), .Z(net_15143) );
SDFFR_X2 inst_2604 ( .D(net_7370), .Q(net_7267), .SI(net_1810), .SE(net_1327), .CK(net_14675), .RN(x6501) );
CLKBUF_X2 inst_18684 ( .A(net_18531), .Z(net_18532) );
CLKBUF_X2 inst_16159 ( .A(net_14426), .Z(net_16007) );
CLKBUF_X2 inst_17776 ( .A(net_17623), .Z(net_17624) );
CLKBUF_X2 inst_15019 ( .A(net_14866), .Z(net_14867) );
NOR4_X2 inst_3248 ( .ZN(net_4383), .A4(net_4320), .A1(net_1467), .A3(net_1431), .A2(net_1104) );
CLKBUF_X2 inst_16961 ( .A(net_16808), .Z(net_16809) );
CLKBUF_X2 inst_18303 ( .A(net_18150), .Z(net_18151) );
CLKBUF_X2 inst_12329 ( .A(net_12137), .Z(net_12177) );
SDFFR_X2 inst_2110 ( .Q(net_7624), .D(net_7624), .SI(net_7623), .SE(net_5750), .CK(net_11127), .RN(x6501) );
CLKBUF_X2 inst_16702 ( .A(net_16549), .Z(net_16550) );
CLKBUF_X2 inst_9774 ( .A(net_9621), .Z(net_9622) );
CLKBUF_X2 inst_13896 ( .A(net_13743), .Z(net_13744) );
DFFR_X1 inst_7463 ( .QN(net_6337), .D(net_4405), .CK(net_17486), .RN(x6501) );
CLKBUF_X2 inst_15051 ( .A(net_14837), .Z(net_14899) );
CLKBUF_X2 inst_18492 ( .A(net_18339), .Z(net_18340) );
CLKBUF_X2 inst_12914 ( .A(net_12314), .Z(net_12762) );
SDFF_X2 inst_2057 ( .SI(net_7923), .Q(net_7923), .D(net_2576), .SE(net_2461), .CK(net_18830) );
CLKBUF_X2 inst_15217 ( .A(net_13304), .Z(net_15065) );
CLKBUF_X2 inst_13408 ( .A(net_10830), .Z(net_13256) );
SDFF_X2 inst_843 ( .SI(net_8654), .Q(net_8654), .D(net_3955), .SE(net_3885), .CK(net_10976) );
CLKBUF_X2 inst_10710 ( .A(net_10557), .Z(net_10558) );
INV_X4 inst_5146 ( .ZN(net_3277), .A(net_3243) );
CLKBUF_X2 inst_14974 ( .A(net_14821), .Z(net_14822) );
SDFF_X2 inst_916 ( .SI(net_8736), .Q(net_8736), .SE(net_6195), .D(net_3950), .CK(net_10507) );
SDFF_X2 inst_1722 ( .Q(net_8185), .D(net_8185), .SI(net_2659), .SE(net_2561), .CK(net_15491) );
INV_X4 inst_5570 ( .A(net_5975), .ZN(net_713) );
CLKBUF_X2 inst_13799 ( .A(net_9380), .Z(net_13647) );
AOI221_X2 inst_8754 ( .ZN(net_5539), .B2(net_5538), .A(net_5276), .C2(net_4388), .C1(net_2624), .B1(net_403) );
DFFR_X2 inst_7300 ( .Q(net_399), .D(net_397), .CK(net_18711), .RN(x6501) );
INV_X2 inst_6409 ( .ZN(net_1066), .A(net_1065) );
NAND4_X2 inst_3665 ( .A4(net_6020), .A1(net_6019), .ZN(net_4600), .A3(net_4102), .A2(net_4101) );
CLKBUF_X2 inst_17433 ( .A(net_17280), .Z(net_17281) );
CLKBUF_X2 inst_16680 ( .A(net_16527), .Z(net_16528) );
CLKBUF_X2 inst_16111 ( .A(net_14040), .Z(net_15959) );
SDFFR_X2 inst_2525 ( .D(net_7372), .SE(net_2387), .SI(net_287), .Q(net_287), .CK(net_16387), .RN(x6501) );
OAI221_X2 inst_2968 ( .C2(net_2650), .B2(net_2649), .ZN(net_2648), .A(net_2646), .C1(net_1273), .B1(net_640) );
CLKBUF_X2 inst_12875 ( .A(net_10509), .Z(net_12723) );
AOI22_X2 inst_7916 ( .A2(net_6426), .A1(net_5654), .ZN(net_4487), .B2(net_4486), .B1(net_568) );
OAI221_X2 inst_2964 ( .ZN(net_3065), .B2(net_3064), .C2(net_3063), .A(net_2882), .C1(net_2350), .B1(net_1447) );
CLKBUF_X2 inst_11760 ( .A(net_9419), .Z(net_11608) );
NAND4_X2 inst_3721 ( .ZN(net_4309), .A1(net_4191), .A2(net_4189), .A4(net_4188), .A3(net_4187) );
SDFFR_X2 inst_2349 ( .SI(net_7369), .SE(net_2732), .D(net_2731), .QN(net_144), .CK(net_16125), .RN(x6501) );
AOI221_X2 inst_8855 ( .B1(net_8882), .C1(net_8327), .B2(net_6252), .ZN(net_6231), .C2(net_4345), .A(net_4244) );
SDFF_X2 inst_646 ( .Q(net_8408), .D(net_8408), .SI(net_3961), .SE(net_3934), .CK(net_10157) );
INV_X4 inst_5076 ( .ZN(net_5849), .A(net_5796) );
HA_X1 inst_6667 ( .S(net_3266), .CO(net_3265), .B(net_3101), .A(x2542) );
NAND2_X4 inst_4032 ( .ZN(net_3086), .A2(net_2903), .A1(net_2902) );
CLKBUF_X2 inst_14310 ( .A(net_14157), .Z(net_14158) );
OAI21_X2 inst_3169 ( .B2(net_1518), .A(net_1515), .ZN(net_1277), .B1(net_862) );
CLKBUF_X2 inst_13278 ( .A(net_13026), .Z(net_13126) );
CLKBUF_X2 inst_9841 ( .A(net_9688), .Z(net_9689) );
INV_X4 inst_5344 ( .ZN(net_1524), .A(net_1114) );
CLKBUF_X2 inst_11119 ( .A(net_10088), .Z(net_10967) );
CLKBUF_X2 inst_14248 ( .A(net_14095), .Z(net_14096) );
CLKBUF_X2 inst_9799 ( .A(net_9646), .Z(net_9647) );
SDFFR_X1 inst_2788 ( .D(net_7393), .Q(net_7290), .SI(net_1960), .SE(net_1327), .CK(net_18334), .RN(x6501) );
INV_X4 inst_6015 ( .A(net_8293), .ZN(net_959) );
CLKBUF_X2 inst_11891 ( .A(net_11738), .Z(net_11739) );
CLKBUF_X2 inst_19191 ( .A(net_19038), .Z(net_19039) );
INV_X2 inst_6565 ( .A(net_6466), .ZN(net_490) );
CLKBUF_X2 inst_10415 ( .A(net_10262), .Z(net_10263) );
CLKBUF_X2 inst_10194 ( .A(net_10041), .Z(net_10042) );
XNOR2_X2 inst_168 ( .ZN(net_1825), .A(net_1544), .B(net_1541) );
AND2_X4 inst_9139 ( .ZN(net_1421), .A2(net_788), .A1(net_179) );
CLKBUF_X2 inst_16173 ( .A(net_16020), .Z(net_16021) );
AOI222_X1 inst_8688 ( .C1(net_6462), .A2(net_3296), .B2(net_3295), .C2(net_3294), .ZN(net_3281), .B1(net_2932), .A1(net_1668) );
SDFF_X2 inst_991 ( .D(net_7329), .SI(net_6637), .Q(net_6637), .SE(net_3123), .CK(net_9525) );
CLKBUF_X2 inst_10642 ( .A(net_10489), .Z(net_10490) );
XNOR2_X2 inst_170 ( .ZN(net_1823), .A(net_1551), .B(net_1548) );
AND2_X2 inst_9160 ( .ZN(net_2808), .A1(net_2807), .A2(net_2806) );
NAND4_X2 inst_3691 ( .ZN(net_4446), .A4(net_4346), .A1(net_3820), .A2(net_3819), .A3(net_3818) );
CLKBUF_X2 inst_17371 ( .A(net_15602), .Z(net_17219) );
CLKBUF_X2 inst_13159 ( .A(net_13006), .Z(net_13007) );
AOI22_X2 inst_7823 ( .B2(net_5463), .A2(net_4881), .ZN(net_4701), .B1(net_440), .A1(net_253) );
SDFF_X2 inst_1857 ( .D(net_7284), .SI(net_6941), .Q(net_6941), .SE(net_6281), .CK(net_16190) );
CLKBUF_X2 inst_11536 ( .A(net_9101), .Z(net_11384) );
SDFF_X2 inst_468 ( .SI(net_8473), .Q(net_8473), .SE(net_3983), .D(net_3953), .CK(net_10287) );
SDFF_X2 inst_1099 ( .D(net_7328), .SI(net_6537), .Q(net_6537), .SE(net_3086), .CK(net_11349) );
CLKBUF_X2 inst_19064 ( .A(net_18911), .Z(net_18912) );
INV_X2 inst_6611 ( .A(net_6200), .ZN(net_6199) );
CLKBUF_X2 inst_17973 ( .A(net_17820), .Z(net_17821) );
NAND2_X2 inst_4428 ( .A1(net_6866), .A2(net_5016), .ZN(net_4999) );
CLKBUF_X2 inst_16805 ( .A(net_16652), .Z(net_16653) );
CLKBUF_X2 inst_14762 ( .A(net_13440), .Z(net_14610) );
NAND2_X2 inst_4889 ( .A2(net_7396), .ZN(net_707), .A1(net_185) );
SDFFR_X2 inst_2190 ( .D(net_2965), .SE(net_2583), .SI(net_2582), .QN(net_289), .CK(net_16426), .RN(x6501) );
SDFF_X2 inst_429 ( .Q(net_8757), .D(net_8757), .SE(net_3982), .SI(net_3944), .CK(net_10852) );
CLKBUF_X2 inst_10298 ( .A(net_10145), .Z(net_10146) );
CLKBUF_X2 inst_18343 ( .A(net_18190), .Z(net_18191) );
CLKBUF_X2 inst_17255 ( .A(net_17102), .Z(net_17103) );
AOI22_X2 inst_7808 ( .A2(net_8228), .B2(net_6144), .ZN(net_4765), .A1(net_4764), .B1(net_4526) );
CLKBUF_X2 inst_18774 ( .A(net_11082), .Z(net_18622) );
INV_X4 inst_5995 ( .A(net_7664), .ZN(net_1549) );
CLKBUF_X2 inst_13824 ( .A(net_9875), .Z(net_13672) );
CLKBUF_X2 inst_13567 ( .A(net_11705), .Z(net_13415) );
CLKBUF_X2 inst_18079 ( .A(net_13891), .Z(net_17927) );
NOR2_X2 inst_3467 ( .ZN(net_2469), .A2(net_2467), .A1(net_790) );
OAI21_X2 inst_3064 ( .B2(net_8220), .B1(net_4850), .ZN(net_4740), .A(net_2625) );
NAND4_X2 inst_3676 ( .A4(net_5992), .A1(net_5991), .ZN(net_4589), .A2(net_4035), .A3(net_4034) );
CLKBUF_X2 inst_15480 ( .A(net_10407), .Z(net_15328) );
AOI22_X2 inst_7948 ( .B1(net_8124), .A1(net_7886), .A2(net_6098), .B2(net_4190), .ZN(net_4178) );
NAND2_X4 inst_4033 ( .ZN(net_3070), .A2(net_2903), .A1(net_2901) );
CLKBUF_X2 inst_18807 ( .A(net_18654), .Z(net_18655) );
CLKBUF_X2 inst_18528 ( .A(net_18375), .Z(net_18376) );
CLKBUF_X2 inst_14210 ( .A(net_14057), .Z(net_14058) );
AOI22_X2 inst_8538 ( .B1(net_6659), .A1(net_6626), .A2(net_6213), .B2(net_6138), .ZN(net_3402) );
INV_X8 inst_5044 ( .ZN(net_6108), .A(net_3560) );
OR2_X2 inst_2899 ( .ZN(net_2466), .A1(net_519), .A2(net_500) );
CLKBUF_X2 inst_15510 ( .A(net_15357), .Z(net_15358) );
CLKBUF_X2 inst_14222 ( .A(net_13736), .Z(net_14070) );
NAND2_X2 inst_4096 ( .ZN(net_5439), .A2(net_5246), .A1(net_5159) );
CLKBUF_X2 inst_10927 ( .A(net_9758), .Z(net_10775) );
DFF_X1 inst_6808 ( .Q(net_8225), .D(net_4420), .CK(net_17225) );
CLKBUF_X2 inst_15323 ( .A(net_15170), .Z(net_15171) );
CLKBUF_X2 inst_12508 ( .A(net_11041), .Z(net_12356) );
SDFF_X2 inst_689 ( .Q(net_8856), .D(net_8856), .SI(net_3938), .SE(net_3936), .CK(net_12437) );
NAND2_X2 inst_4453 ( .ZN(net_4963), .A2(net_4962), .A1(net_3254) );
SDFFR_X1 inst_2689 ( .SI(net_7552), .SE(net_5043), .CK(net_12747), .RN(x6501), .Q(x3891), .D(x3891) );
CLKBUF_X2 inst_16306 ( .A(net_15794), .Z(net_16154) );
CLKBUF_X2 inst_16123 ( .A(net_15970), .Z(net_15971) );
CLKBUF_X2 inst_9622 ( .A(net_9469), .Z(net_9470) );
CLKBUF_X2 inst_12630 ( .A(net_12477), .Z(net_12478) );
CLKBUF_X2 inst_18499 ( .A(net_18346), .Z(net_18347) );
INV_X2 inst_6272 ( .A(net_6328), .ZN(net_4405) );
CLKBUF_X2 inst_17532 ( .A(net_17122), .Z(net_17380) );
CLKBUF_X2 inst_13587 ( .A(net_13434), .Z(net_13435) );
AOI222_X1 inst_8685 ( .B1(net_6484), .A2(net_3296), .B2(net_3295), .C2(net_3294), .ZN(net_3287), .C1(net_3286), .A1(net_1215) );
SDFF_X2 inst_1615 ( .Q(net_8156), .D(net_8156), .SI(net_2584), .SE(net_2538), .CK(net_18859) );
CLKBUF_X2 inst_16718 ( .A(net_12603), .Z(net_16566) );
AND2_X4 inst_9148 ( .A2(net_7483), .A1(net_7481), .ZN(net_1657) );
CLKBUF_X2 inst_11434 ( .A(net_9190), .Z(net_11282) );
DFFR_X1 inst_7503 ( .Q(net_7264), .D(net_1878), .CK(net_17485), .RN(x6501) );
CLKBUF_X2 inst_12406 ( .A(net_10052), .Z(net_12254) );
CLKBUF_X2 inst_13760 ( .A(net_13607), .Z(net_13608) );
AOI22_X2 inst_8313 ( .B1(net_8743), .A1(net_8373), .A2(net_3867), .B2(net_3866), .ZN(net_3732) );
SDFFR_X2 inst_2145 ( .SI(net_7172), .Q(net_7172), .SE(net_3586), .D(net_3026), .CK(net_15153), .RN(x6501) );
CLKBUF_X2 inst_17890 ( .A(net_17737), .Z(net_17738) );
SDFF_X2 inst_709 ( .SI(net_8617), .Q(net_8617), .SE(net_3984), .D(net_3955), .CK(net_13242) );
SDFFR_X2 inst_2375 ( .SE(net_2260), .Q(net_322), .D(net_322), .CK(net_10432), .RN(x6501), .SI(x3028) );
INV_X4 inst_5725 ( .A(net_7262), .ZN(net_566) );
CLKBUF_X2 inst_18431 ( .A(net_13146), .Z(net_18279) );
CLKBUF_X2 inst_13400 ( .A(net_12097), .Z(net_13248) );
CLKBUF_X2 inst_12080 ( .A(net_11927), .Z(net_11928) );
CLKBUF_X2 inst_9956 ( .A(net_9803), .Z(net_9804) );
CLKBUF_X2 inst_12517 ( .A(net_12364), .Z(net_12365) );
CLKBUF_X2 inst_12331 ( .A(net_9369), .Z(net_12179) );
CLKBUF_X2 inst_12106 ( .A(net_10140), .Z(net_11954) );
DFFR_X1 inst_7389 ( .D(net_5857), .CK(net_14060), .RN(x6501), .Q(x406) );
NAND2_X2 inst_4610 ( .A2(net_6144), .ZN(net_2621), .A1(net_2620) );
CLKBUF_X2 inst_13350 ( .A(net_13197), .Z(net_13198) );
NAND2_X2 inst_4403 ( .A1(net_7047), .A2(net_5162), .ZN(net_5054) );
CLKBUF_X2 inst_19076 ( .A(net_16542), .Z(net_18924) );
CLKBUF_X2 inst_14589 ( .A(net_14277), .Z(net_14437) );
CLKBUF_X2 inst_11432 ( .A(net_11279), .Z(net_11280) );
CLKBUF_X2 inst_9885 ( .A(net_9732), .Z(net_9733) );
OAI22_X2 inst_2935 ( .B2(net_2282), .A2(net_2146), .ZN(net_2095), .B1(net_2031), .A1(net_1428) );
NOR2_X2 inst_3369 ( .ZN(net_5556), .A1(net_5352), .A2(net_5351) );
CLKBUF_X2 inst_13612 ( .A(net_11408), .Z(net_13460) );
CLKBUF_X2 inst_17545 ( .A(net_13265), .Z(net_17393) );
CLKBUF_X2 inst_16507 ( .A(net_14855), .Z(net_16355) );
CLKBUF_X2 inst_10924 ( .A(net_10771), .Z(net_10772) );
CLKBUF_X2 inst_14444 ( .A(net_14291), .Z(net_14292) );
AND2_X2 inst_9202 ( .A1(net_8214), .ZN(net_1455), .A2(net_743) );
CLKBUF_X2 inst_10179 ( .A(net_10026), .Z(net_10027) );
SDFF_X2 inst_415 ( .SI(net_8329), .Q(net_8329), .SE(net_3978), .D(net_3950), .CK(net_13290) );
CLKBUF_X2 inst_10592 ( .A(net_10119), .Z(net_10440) );
CLKBUF_X2 inst_17508 ( .A(net_9912), .Z(net_17356) );
CLKBUF_X2 inst_12005 ( .A(net_10574), .Z(net_11853) );
AOI22_X2 inst_7866 ( .B2(net_4881), .A2(net_4809), .ZN(net_4575), .A1(net_349), .B1(net_255) );
DFFR_X2 inst_7291 ( .D(net_394), .QN(net_391), .CK(net_13863), .RN(x6501) );
CLKBUF_X2 inst_17348 ( .A(net_17195), .Z(net_17196) );
CLKBUF_X2 inst_15772 ( .A(net_15226), .Z(net_15620) );
AND2_X4 inst_9074 ( .ZN(net_3378), .A1(net_3180), .A2(net_3179) );
INV_X2 inst_6278 ( .ZN(net_4270), .A(net_4225) );
CLKBUF_X2 inst_16601 ( .A(net_16448), .Z(net_16449) );
CLKBUF_X2 inst_15494 ( .A(net_15341), .Z(net_15342) );
CLKBUF_X2 inst_10869 ( .A(net_10716), .Z(net_10717) );
CLKBUF_X2 inst_14185 ( .A(net_9270), .Z(net_14033) );
CLKBUF_X2 inst_10408 ( .A(net_9970), .Z(net_10256) );
SDFF_X2 inst_1561 ( .Q(net_7898), .D(net_7898), .SI(net_2717), .SE(net_2543), .CK(net_14177) );
SDFFR_X2 inst_2104 ( .SE(net_5921), .SI(net_5920), .Q(net_388), .D(net_388), .CK(net_17555), .RN(x6501) );
CLKBUF_X2 inst_12190 ( .A(net_12037), .Z(net_12038) );
CLKBUF_X2 inst_12437 ( .A(net_12284), .Z(net_12285) );
CLKBUF_X2 inst_9530 ( .A(net_9235), .Z(net_9378) );
SDFFR_X2 inst_2573 ( .SI(net_6833), .Q(net_6833), .D(net_6830), .SE(net_2146), .CK(net_18688), .RN(x6501) );
CLKBUF_X2 inst_16701 ( .A(net_16548), .Z(net_16549) );
AOI221_X2 inst_8762 ( .C2(net_6130), .B2(net_5535), .ZN(net_5470), .A(net_4946), .C1(net_1397), .B1(net_462) );
CLKBUF_X1 inst_7733 ( .A(x192486), .Z(x4227) );
INV_X2 inst_6233 ( .ZN(net_5477), .A(net_5294) );
CLKBUF_X2 inst_14760 ( .A(net_14607), .Z(net_14608) );
CLKBUF_X2 inst_14564 ( .A(net_12010), .Z(net_14412) );
SDFFS_X2 inst_2096 ( .Q(net_7522), .D(net_7522), .SI(net_2068), .SE(net_1136), .CK(net_16246), .SN(x6501) );
CLKBUF_X2 inst_10169 ( .A(net_10016), .Z(net_10017) );
SDFF_X2 inst_552 ( .Q(net_8698), .D(net_8698), .SI(net_3951), .SE(net_3935), .CK(net_12890) );
NAND2_X2 inst_4793 ( .ZN(net_1868), .A1(net_1500), .A2(net_1109) );
CLKBUF_X2 inst_18394 ( .A(net_18241), .Z(net_18242) );
MUX2_X2 inst_4997 ( .A(net_9029), .Z(net_3959), .B(net_2921), .S(net_622) );
CLKBUF_X2 inst_12483 ( .A(net_10279), .Z(net_12331) );
SDFF_X2 inst_1564 ( .Q(net_8013), .D(net_8013), .SI(net_2655), .SE(net_2545), .CK(net_15437) );
DFFR_X2 inst_6985 ( .D(net_5892), .CK(net_11441), .RN(x6501), .Q(x2308) );
CLKBUF_X2 inst_10995 ( .A(net_10018), .Z(net_10843) );
CLKBUF_X2 inst_18256 ( .A(net_10678), .Z(net_18104) );
INV_X2 inst_6477 ( .ZN(net_815), .A(net_215) );
AOI22_X2 inst_8064 ( .B1(net_8072), .A1(net_7868), .B2(net_6107), .ZN(net_6024), .A2(net_4400) );
CLKBUF_X2 inst_15260 ( .A(net_15107), .Z(net_15108) );
CLKBUF_X2 inst_9492 ( .A(net_9172), .Z(net_9340) );
SDFF_X2 inst_356 ( .Q(net_8767), .D(net_8767), .SE(net_3982), .SI(net_3975), .CK(net_12572) );
CLKBUF_X2 inst_9311 ( .A(net_9058), .Z(net_9159) );
CLKBUF_X2 inst_17627 ( .A(net_11838), .Z(net_17475) );
INV_X4 inst_5587 ( .A(net_7500), .ZN(net_3205) );
CLKBUF_X2 inst_10735 ( .A(net_10582), .Z(net_10583) );
CLKBUF_X2 inst_16696 ( .A(net_16543), .Z(net_16544) );
DFFS_X2 inst_6884 ( .QN(net_6155), .D(net_3117), .CK(net_18474), .SN(x6501) );
CLKBUF_X2 inst_9267 ( .A(net_9114), .Z(net_9115) );
AND2_X4 inst_9105 ( .A2(net_2299), .ZN(net_2267), .A1(net_1455) );
NAND2_X2 inst_4286 ( .A1(net_7008), .A2(net_5249), .ZN(net_5174) );
CLKBUF_X2 inst_16004 ( .A(net_15851), .Z(net_15852) );
SDFF_X2 inst_1935 ( .SI(net_8065), .Q(net_8065), .D(net_2713), .SE(net_2508), .CK(net_16462) );
INV_X4 inst_6032 ( .A(net_7565), .ZN(net_503) );
CLKBUF_X2 inst_9332 ( .A(net_9148), .Z(net_9180) );
CLKBUF_X2 inst_14949 ( .A(net_14796), .Z(net_14797) );
AOI222_X1 inst_8678 ( .ZN(net_3298), .A2(net_3296), .B2(net_3295), .C2(net_3294), .C1(net_3292), .B1(net_2770), .A1(net_1233) );
CLKBUF_X2 inst_19133 ( .A(net_18980), .Z(net_18981) );
AOI22_X2 inst_8235 ( .B1(net_8686), .A1(net_8649), .B2(net_6109), .A2(net_3857), .ZN(net_3802) );
CLKBUF_X2 inst_15927 ( .A(net_13378), .Z(net_15775) );
CLKBUF_X2 inst_13884 ( .A(net_13731), .Z(net_13732) );
SDFFR_X2 inst_2140 ( .SI(net_7180), .Q(net_7180), .D(net_6431), .SE(net_4362), .CK(net_16431), .RN(x6501) );
CLKBUF_X2 inst_14501 ( .A(net_10270), .Z(net_14349) );
CLKBUF_X2 inst_9641 ( .A(net_9488), .Z(net_9489) );
CLKBUF_X2 inst_11386 ( .A(net_11233), .Z(net_11234) );
CLKBUF_X2 inst_9499 ( .A(net_9346), .Z(net_9347) );
CLKBUF_X2 inst_15648 ( .A(net_15495), .Z(net_15496) );
CLKBUF_X2 inst_13120 ( .A(net_12967), .Z(net_12968) );
CLKBUF_X2 inst_19130 ( .A(net_18977), .Z(net_18978) );
SDFF_X2 inst_1559 ( .Q(net_7879), .D(net_7879), .SI(net_2659), .SE(net_2543), .CK(net_15525) );
AOI221_X2 inst_8830 ( .B1(net_8063), .C1(net_7859), .B2(net_6107), .ZN(net_6009), .C2(net_4400), .A(net_4300) );
DFF_X1 inst_6752 ( .Q(net_6762), .D(net_5614), .CK(net_10493) );
SDFF_X2 inst_927 ( .SI(net_8728), .Q(net_8728), .SE(net_6195), .D(net_3955), .CK(net_13230) );
CLKBUF_X2 inst_13304 ( .A(net_9683), .Z(net_13152) );
DFFR_X1 inst_7420 ( .D(net_5468), .CK(net_16615), .RN(x6501), .Q(x649) );
CLKBUF_X2 inst_13258 ( .A(net_13105), .Z(net_13106) );
XOR2_X1 inst_73 ( .B(net_4465), .Z(net_3384), .A(net_3222) );
SDFF_X2 inst_1488 ( .SI(net_7295), .Q(net_7072), .D(net_7072), .SE(net_6280), .CK(net_15450) );
SDFF_X2 inst_1719 ( .Q(net_8000), .D(net_8000), .SI(net_2717), .SE(net_2542), .CK(net_14398) );
NAND2_X2 inst_4690 ( .ZN(net_1991), .A1(net_1928), .A2(net_1769) );
CLKBUF_X2 inst_9236 ( .A(net_9083), .Z(net_9084) );
SDFF_X2 inst_890 ( .Q(net_8582), .D(net_8582), .SI(net_3975), .SE(net_3878), .CK(net_12488) );
CLKBUF_X2 inst_12510 ( .A(net_9368), .Z(net_12358) );
CLKBUF_X2 inst_12352 ( .A(net_12199), .Z(net_12200) );
SDFF_X2 inst_1851 ( .D(net_7273), .SI(net_6930), .Q(net_6930), .SE(net_6281), .CK(net_14107) );
INV_X4 inst_5911 ( .ZN(net_1817), .A(net_270) );
CLKBUF_X2 inst_12896 ( .A(net_12743), .Z(net_12744) );
NAND2_X2 inst_4514 ( .ZN(net_4315), .A2(net_4272), .A1(net_2846) );
CLKBUF_X2 inst_18842 ( .A(net_18689), .Z(net_18690) );
DFFS_X2 inst_6903 ( .Q(net_7166), .D(net_2095), .CK(net_18703), .SN(x6501) );
SDFF_X2 inst_1168 ( .D(net_7328), .SI(net_6504), .Q(net_6504), .SE(net_3071), .CK(net_11749) );
CLKBUF_X2 inst_12963 ( .A(net_12810), .Z(net_12811) );
CLKBUF_X2 inst_17808 ( .A(net_14203), .Z(net_17656) );
CLKBUF_X2 inst_15395 ( .A(net_13518), .Z(net_15243) );
CLKBUF_X2 inst_15092 ( .A(net_14939), .Z(net_14940) );
NAND2_X2 inst_4363 ( .A1(net_7111), .A2(net_5164), .ZN(net_5094) );
SDFF_X2 inst_1161 ( .SI(net_7314), .Q(net_6589), .D(net_6589), .SE(net_3069), .CK(net_9901) );
NOR2_X2 inst_3362 ( .ZN(net_5563), .A1(net_5380), .A2(net_5379) );
CLKBUF_X2 inst_17743 ( .A(net_17590), .Z(net_17591) );
CLKBUF_X2 inst_17308 ( .A(net_17155), .Z(net_17156) );
CLKBUF_X2 inst_17177 ( .A(net_17024), .Z(net_17025) );
CLKBUF_X2 inst_15667 ( .A(net_15514), .Z(net_15515) );
CLKBUF_X2 inst_17521 ( .A(net_17368), .Z(net_17369) );
CLKBUF_X2 inst_17897 ( .A(net_9461), .Z(net_17745) );
CLKBUF_X2 inst_14096 ( .A(net_10027), .Z(net_13944) );
CLKBUF_X2 inst_18062 ( .A(net_17909), .Z(net_17910) );
CLKBUF_X2 inst_16739 ( .A(net_16586), .Z(net_16587) );
CLKBUF_X2 inst_10703 ( .A(net_10550), .Z(net_10551) );
SDFFR_X2 inst_2388 ( .SE(net_2260), .Q(net_367), .D(net_367), .CK(net_9288), .RN(x6501), .SI(x1745) );
CLKBUF_X2 inst_15984 ( .A(net_15831), .Z(net_15832) );
INV_X4 inst_5633 ( .A(net_7367), .ZN(net_1877) );
NAND2_X2 inst_4309 ( .A1(net_7095), .A2(net_5164), .ZN(net_5148) );
CLKBUF_X2 inst_11642 ( .A(net_11489), .Z(net_11490) );
SDFFR_X2 inst_2634 ( .Q(net_7367), .D(net_7367), .SE(net_1136), .CK(net_18605), .RN(x6501), .SI(x4851) );
NAND4_X2 inst_3711 ( .ZN(net_4426), .A4(net_4333), .A1(net_3694), .A2(net_3693), .A3(net_3692) );
CLKBUF_X2 inst_16812 ( .A(net_16659), .Z(net_16660) );
CLKBUF_X2 inst_16408 ( .A(net_16255), .Z(net_16256) );
CLKBUF_X2 inst_17178 ( .A(net_17025), .Z(net_17026) );
DFFR_X1 inst_7568 ( .D(net_7626), .QN(net_7625), .CK(net_11261), .RN(x6501) );
SDFF_X2 inst_650 ( .Q(net_8421), .D(net_8421), .SI(net_3966), .SE(net_3934), .CK(net_10001) );
XNOR2_X2 inst_289 ( .B(net_1023), .ZN(net_1003), .A(net_535) );
AOI222_X1 inst_8674 ( .C1(net_7512), .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3385), .A2(net_3197), .B1(net_3135) );
CLKBUF_X2 inst_12467 ( .A(net_12314), .Z(net_12315) );
AOI222_X1 inst_8701 ( .A2(net_8251), .C2(net_6116), .A1(net_4800), .B2(net_4799), .ZN(net_2837), .B1(net_2836), .C1(net_2569) );
AOI222_X1 inst_8643 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3930), .B1(net_2463), .C1(net_2462), .A1(x13843) );
SDFF_X2 inst_679 ( .Q(net_8699), .D(net_8699), .SI(net_3950), .SE(net_3935), .CK(net_12607) );
CLKBUF_X2 inst_17472 ( .A(net_17319), .Z(net_17320) );
INV_X4 inst_5627 ( .A(net_8934), .ZN(net_2632) );
CLKBUF_X2 inst_16666 ( .A(net_16513), .Z(net_16514) );
CLKBUF_X2 inst_12532 ( .A(net_12379), .Z(net_12380) );
NOR2_X2 inst_3364 ( .ZN(net_5561), .A1(net_5372), .A2(net_5371) );
SDFF_X2 inst_1351 ( .Q(net_8198), .D(net_8198), .SI(net_2590), .SE(net_2561), .CK(net_18805) );
CLKBUF_X2 inst_10443 ( .A(net_9884), .Z(net_10291) );
XOR2_X2 inst_44 ( .A(net_7590), .Z(net_1038), .B(net_1037) );
NAND2_X2 inst_4433 ( .A1(net_6870), .A2(net_5016), .ZN(net_4994) );
CLKBUF_X2 inst_16501 ( .A(net_16348), .Z(net_16349) );
CLKBUF_X2 inst_13994 ( .A(net_9591), .Z(net_13842) );
CLKBUF_X2 inst_12805 ( .A(net_12193), .Z(net_12653) );
SDFF_X2 inst_435 ( .Q(net_8763), .D(net_8763), .SE(net_3982), .SI(net_3963), .CK(net_10942) );
CLKBUF_X2 inst_11563 ( .A(net_11410), .Z(net_11411) );
CLKBUF_X2 inst_10791 ( .A(net_10638), .Z(net_10639) );
CLKBUF_X2 inst_10305 ( .A(net_9758), .Z(net_10153) );
CLKBUF_X2 inst_13474 ( .A(net_13321), .Z(net_13322) );
NAND4_X2 inst_3787 ( .A3(net_6071), .A1(net_6070), .ZN(net_4234), .A2(net_3657), .A4(net_3656) );
MUX2_X2 inst_4982 ( .A(net_9043), .Z(net_3953), .B(net_652), .S(net_622) );
CLKBUF_X2 inst_13633 ( .A(net_9237), .Z(net_13481) );
SDFF_X2 inst_1923 ( .D(net_7287), .SI(net_7024), .Q(net_7024), .SE(net_6277), .CK(net_18753) );
SDFFR_X1 inst_2748 ( .SI(net_9036), .Q(net_9036), .D(net_7465), .SE(net_3208), .CK(net_10646), .RN(x6501) );
OAI21_X2 inst_3013 ( .ZN(net_5527), .A(net_5271), .B2(net_5270), .B1(x1130) );
AND2_X2 inst_9201 ( .A2(net_1619), .ZN(net_1279), .A1(net_881) );
NAND2_X2 inst_4744 ( .ZN(net_2660), .A2(net_1586), .A1(net_1126) );
INV_X4 inst_5087 ( .ZN(net_5726), .A(net_5699) );
AND2_X4 inst_9130 ( .ZN(net_1409), .A2(net_851), .A1(net_184) );
DFFR_X1 inst_7563 ( .Q(net_398), .D(net_269), .CK(net_11627), .RN(x6501) );
CLKBUF_X2 inst_14656 ( .A(net_14503), .Z(net_14504) );
CLKBUF_X2 inst_11127 ( .A(net_10974), .Z(net_10975) );
CLKBUF_X2 inst_13931 ( .A(net_11348), .Z(net_13779) );
SDFFR_X1 inst_2734 ( .SI(net_9048), .Q(net_9048), .SE(net_3208), .D(net_3129), .CK(net_10655), .RN(x6501) );
MUX2_X2 inst_4920 ( .S(net_6272), .Z(net_4623), .A(net_4622), .B(net_4621) );
CLKBUF_X2 inst_14956 ( .A(net_9177), .Z(net_14804) );
CLKBUF_X2 inst_18959 ( .A(net_18806), .Z(net_18807) );
CLKBUF_X2 inst_11608 ( .A(net_11455), .Z(net_11456) );
INV_X2 inst_6518 ( .ZN(net_886), .A(net_213) );
SDFF_X2 inst_855 ( .SI(net_8635), .Q(net_8635), .D(net_3965), .SE(net_3885), .CK(net_12414) );
SDFF_X2 inst_2039 ( .SI(net_7785), .Q(net_7785), .D(net_2720), .SE(net_2459), .CK(net_15472) );
CLKBUF_X2 inst_15241 ( .A(net_15040), .Z(net_15089) );
NOR4_X2 inst_3233 ( .ZN(net_2023), .A2(net_1735), .A1(net_1420), .A3(net_1404), .A4(net_1402) );
CLKBUF_X2 inst_15226 ( .A(net_15073), .Z(net_15074) );
INV_X4 inst_5866 ( .A(net_9056), .ZN(net_2913) );
INV_X4 inst_5466 ( .ZN(net_758), .A(net_757) );
CLKBUF_X2 inst_10160 ( .A(net_10007), .Z(net_10008) );
NAND2_X2 inst_4295 ( .A1(net_7050), .ZN(net_5163), .A2(net_5162) );
SDFF_X2 inst_518 ( .Q(net_8872), .D(net_8872), .SI(net_3957), .SE(net_3936), .CK(net_13263) );
CLKBUF_X2 inst_19196 ( .A(net_19043), .Z(net_19044) );
INV_X4 inst_5894 ( .ZN(net_3542), .A(net_476) );
AOI22_X2 inst_8242 ( .B1(net_8668), .A1(net_8631), .B2(net_6109), .A2(net_3857), .ZN(net_3795) );
NAND4_X2 inst_3863 ( .ZN(net_1345), .A3(x2594), .A4(x2542), .A1(x2494), .A2(x2451) );
SDFFR_X2 inst_2345 ( .D(net_7367), .SE(net_2734), .SI(net_273), .Q(net_273), .CK(net_13684), .RN(x6501) );
CLKBUF_X2 inst_12157 ( .A(net_12004), .Z(net_12005) );
CLKBUF_X2 inst_18081 ( .A(net_17928), .Z(net_17929) );
INV_X2 inst_6538 ( .A(net_5945), .ZN(x1195) );
NOR2_X2 inst_3602 ( .A2(net_7619), .ZN(net_3251), .A1(net_492) );
CLKBUF_X2 inst_9614 ( .A(net_9461), .Z(net_9462) );
CLKBUF_X2 inst_15967 ( .A(net_15814), .Z(net_15815) );
CLKBUF_X2 inst_14291 ( .A(net_14138), .Z(net_14139) );
DFFR_X1 inst_7582 ( .D(net_6414), .QN(net_6413), .CK(net_15211), .RN(x6501) );
INV_X4 inst_5260 ( .ZN(net_2047), .A(net_1876) );
CLKBUF_X2 inst_12637 ( .A(net_12484), .Z(net_12485) );
CLKBUF_X2 inst_11815 ( .A(net_11662), .Z(net_11663) );
CLKBUF_X2 inst_17291 ( .A(net_10326), .Z(net_17139) );
CLKBUF_X2 inst_12336 ( .A(net_12183), .Z(net_12184) );
INV_X4 inst_5190 ( .ZN(net_2933), .A(net_2897) );
SDFF_X2 inst_1354 ( .Q(net_8193), .D(net_8193), .SI(net_2720), .SE(net_2561), .CK(net_18071) );
SDFF_X2 inst_970 ( .SI(net_7331), .Q(net_6738), .D(net_6738), .SE(net_3124), .CK(net_9080) );
CLKBUF_X2 inst_18088 ( .A(net_11399), .Z(net_17936) );
DFF_X1 inst_6731 ( .Q(net_6776), .D(net_5638), .CK(net_9209) );
SDFF_X2 inst_1278 ( .Q(net_7836), .D(net_7836), .SE(net_2730), .SI(net_2704), .CK(net_17026) );
NAND4_X2 inst_3763 ( .ZN(net_4258), .A1(net_3811), .A2(net_3810), .A3(net_3809), .A4(net_3808) );
CLKBUF_X2 inst_10136 ( .A(net_9291), .Z(net_9984) );
SDFF_X2 inst_749 ( .Q(net_8788), .D(net_8788), .SI(net_3960), .SE(net_3879), .CK(net_12256) );
CLKBUF_X2 inst_15159 ( .A(net_10027), .Z(net_15007) );
CLKBUF_X2 inst_11975 ( .A(net_11822), .Z(net_11823) );
SDFF_X2 inst_1030 ( .D(net_7318), .SI(net_6626), .Q(net_6626), .SE(net_3123), .CK(net_12108) );
SDFFR_X1 inst_2649 ( .D(net_6772), .SE(net_4506), .CK(net_9237), .RN(x6501), .SI(x1721), .Q(x1721) );
CLKBUF_X2 inst_11441 ( .A(net_11288), .Z(net_11289) );
NAND4_X2 inst_3828 ( .ZN(net_2765), .A4(net_2336), .A2(net_2276), .A3(net_2110), .A1(net_1782) );
INV_X4 inst_5841 ( .A(net_6392), .ZN(net_1762) );
DFFS_X2 inst_6898 ( .Q(net_8953), .D(net_2572), .CK(net_17232), .SN(x6501) );
CLKBUF_X2 inst_17006 ( .A(net_13591), .Z(net_16854) );
SDFF_X2 inst_1006 ( .D(net_7317), .SI(net_6625), .Q(net_6625), .SE(net_3123), .CK(net_9871) );
SDFF_X2 inst_1985 ( .D(net_7290), .SI(net_7027), .Q(net_7027), .SE(net_6277), .CK(net_15303) );
DFFR_X2 inst_7311 ( .D(net_292), .QN(net_151), .CK(net_11140), .RN(x6501) );
CLKBUF_X2 inst_17981 ( .A(net_12088), .Z(net_17829) );
CLKBUF_X2 inst_14878 ( .A(net_14341), .Z(net_14726) );
CLKBUF_X2 inst_13519 ( .A(net_12195), .Z(net_13367) );
CLKBUF_X2 inst_10473 ( .A(net_10320), .Z(net_10321) );
CLKBUF_X2 inst_9817 ( .A(net_9450), .Z(net_9665) );
INV_X4 inst_5134 ( .ZN(net_4272), .A(net_4216) );
DFFR_X2 inst_7180 ( .QN(net_8951), .D(net_2469), .CK(net_17236), .RN(x6501) );
AOI222_X1 inst_8691 ( .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3237), .C1(net_3236), .B1(net_3139), .A2(net_3041) );
NAND2_X2 inst_4753 ( .ZN(net_2720), .A1(net_1745), .A2(net_1586) );
CLKBUF_X2 inst_10960 ( .A(net_10807), .Z(net_10808) );
CLKBUF_X2 inst_16168 ( .A(net_16015), .Z(net_16016) );
CLKBUF_X2 inst_11885 ( .A(net_10898), .Z(net_11733) );
CLKBUF_X2 inst_10082 ( .A(net_9387), .Z(net_9930) );
CLKBUF_X2 inst_11957 ( .A(net_10813), .Z(net_11805) );
MUX2_X2 inst_4947 ( .A(net_7396), .Z(net_2379), .S(net_2378), .B(net_905) );
AOI21_X2 inst_8915 ( .B2(net_5784), .ZN(net_5722), .A(net_5721), .B1(net_2736) );
CLKBUF_X2 inst_11671 ( .A(net_11468), .Z(net_11519) );
CLKBUF_X2 inst_15986 ( .A(net_15833), .Z(net_15834) );
CLKBUF_X2 inst_18456 ( .A(net_18303), .Z(net_18304) );
CLKBUF_X2 inst_18208 ( .A(net_18055), .Z(net_18056) );
INV_X4 inst_5783 ( .A(net_6353), .ZN(net_548) );
CLKBUF_X2 inst_16413 ( .A(net_16260), .Z(net_16261) );
CLKBUF_X2 inst_15701 ( .A(net_15548), .Z(net_15549) );
INV_X2 inst_6457 ( .A(net_6486), .ZN(net_585) );
CLKBUF_X2 inst_9898 ( .A(net_9745), .Z(net_9746) );
NAND2_X2 inst_4184 ( .ZN(net_5318), .A1(net_5187), .A2(net_4986) );
INV_X2 inst_6531 ( .A(net_7524), .ZN(net_1083) );
CLKBUF_X2 inst_11517 ( .A(net_9399), .Z(net_11365) );
NOR4_X2 inst_3238 ( .A1(net_1976), .ZN(net_1781), .A4(net_1701), .A2(net_1585), .A3(net_1309) );
OR2_X4 inst_2854 ( .ZN(net_3161), .A2(net_882), .A1(net_880) );
OAI21_X2 inst_3030 ( .B1(net_4954), .ZN(net_4931), .B2(net_4853), .A(net_4717) );
SDFFR_X2 inst_2230 ( .Q(net_7468), .D(net_7468), .SE(net_2863), .CK(net_12170), .SI(x13447), .RN(x6501) );
INV_X4 inst_5630 ( .A(net_8937), .ZN(net_4540) );
CLKBUF_X2 inst_13028 ( .A(net_12875), .Z(net_12876) );
CLKBUF_X2 inst_18621 ( .A(net_18468), .Z(net_18469) );
CLKBUF_X2 inst_17512 ( .A(net_17359), .Z(net_17360) );
CLKBUF_X2 inst_10511 ( .A(net_10358), .Z(net_10359) );
CLKBUF_X2 inst_13820 ( .A(net_13667), .Z(net_13668) );
CLKBUF_X2 inst_10481 ( .A(net_10328), .Z(net_10329) );
CLKBUF_X2 inst_14964 ( .A(net_13706), .Z(net_14812) );
CLKBUF_X2 inst_18153 ( .A(net_18000), .Z(net_18001) );
CLKBUF_X2 inst_14174 ( .A(net_14021), .Z(net_14022) );
NAND2_X2 inst_4477 ( .ZN(net_4507), .A2(net_4388), .A1(net_2610) );
SDFFR_X2 inst_2391 ( .SE(net_2260), .Q(net_354), .D(net_354), .CK(net_10415), .RN(x6501), .SI(x2133) );
CLKBUF_X2 inst_17588 ( .A(net_10463), .Z(net_17436) );
CLKBUF_X2 inst_14837 ( .A(net_11170), .Z(net_14685) );
SDFFR_X2 inst_2239 ( .Q(net_7454), .D(net_7454), .SE(net_2863), .CK(net_12917), .SI(x13547), .RN(x6501) );
CLKBUF_X2 inst_15601 ( .A(net_15448), .Z(net_15449) );
CLKBUF_X2 inst_10027 ( .A(net_9874), .Z(net_9875) );
INV_X2 inst_6335 ( .A(net_3928), .ZN(net_2887) );
SDFF_X2 inst_1639 ( .Q(net_8155), .D(net_8155), .SI(net_2573), .SE(net_2538), .CK(net_15508) );
CLKBUF_X2 inst_13645 ( .A(net_13492), .Z(net_13493) );
CLKBUF_X2 inst_11468 ( .A(net_11315), .Z(net_11316) );
CLKBUF_X2 inst_10717 ( .A(net_9692), .Z(net_10565) );
CLKBUF_X2 inst_15443 ( .A(net_14994), .Z(net_15291) );
CLKBUF_X2 inst_14743 ( .A(net_14590), .Z(net_14591) );
INV_X4 inst_5155 ( .ZN(net_3260), .A(net_3220) );
CLKBUF_X2 inst_10365 ( .A(net_10212), .Z(net_10213) );
CLKBUF_X2 inst_11071 ( .A(net_10918), .Z(net_10919) );
CLKBUF_X2 inst_9756 ( .A(net_9603), .Z(net_9604) );
DFFR_X1 inst_7403 ( .D(net_5728), .CK(net_13904), .RN(x6501), .Q(x577) );
XNOR2_X2 inst_155 ( .A(net_2146), .ZN(net_2016), .B(net_2015) );
NAND2_X2 inst_4858 ( .ZN(net_1417), .A2(net_886), .A1(net_169) );
CLKBUF_X2 inst_10170 ( .A(net_10017), .Z(net_10018) );
INV_X4 inst_6043 ( .A(net_6287), .ZN(net_2677) );
INV_X4 inst_5309 ( .ZN(net_1700), .A(net_1477) );
XOR2_X2 inst_55 ( .A(net_3170), .Z(net_982), .B(net_559) );
SDFFR_X2 inst_2280 ( .SI(net_7393), .SE(net_2789), .Q(net_252), .D(net_252), .CK(net_17759), .RN(x6501) );
CLKBUF_X2 inst_9872 ( .A(net_9542), .Z(net_9720) );
DFFR_X2 inst_7097 ( .Q(net_6462), .D(net_3339), .CK(net_15105), .RN(x6501) );
NAND2_X2 inst_4127 ( .ZN(net_5397), .A1(net_5225), .A2(net_5005) );
CLKBUF_X2 inst_17786 ( .A(net_17633), .Z(net_17634) );
CLKBUF_X2 inst_17440 ( .A(net_17287), .Z(net_17288) );
CLKBUF_X2 inst_11634 ( .A(net_9500), .Z(net_11482) );
XNOR2_X2 inst_323 ( .B(net_1007), .ZN(net_937), .A(net_936) );
SDFF_X2 inst_1494 ( .SI(net_7850), .Q(net_7850), .D(net_2584), .SE(net_2558), .CK(net_18866) );
CLKBUF_X2 inst_17792 ( .A(net_17639), .Z(net_17640) );
NOR2_X2 inst_3525 ( .A1(net_4320), .A2(net_3262), .ZN(net_1708) );
CLKBUF_X2 inst_12734 ( .A(net_12581), .Z(net_12582) );
CLKBUF_X2 inst_10479 ( .A(net_10326), .Z(net_10327) );
NOR2_X2 inst_3449 ( .A1(net_3023), .ZN(net_2982), .A2(net_2879) );
CLKBUF_X2 inst_18236 ( .A(net_17817), .Z(net_18084) );
CLKBUF_X2 inst_17748 ( .A(net_17595), .Z(net_17596) );
CLKBUF_X2 inst_17332 ( .A(net_11756), .Z(net_17180) );
SDFF_X2 inst_1340 ( .Q(net_8194), .D(net_8194), .SI(net_2589), .SE(net_2561), .CK(net_15613) );
SDFF_X2 inst_1481 ( .SI(net_7266), .Q(net_7083), .D(net_7083), .SE(net_6278), .CK(net_14363) );
CLKBUF_X2 inst_14275 ( .A(net_14122), .Z(net_14123) );
CLKBUF_X2 inst_18326 ( .A(net_18173), .Z(net_18174) );
CLKBUF_X2 inst_18563 ( .A(net_18410), .Z(net_18411) );
CLKBUF_X2 inst_14785 ( .A(net_13624), .Z(net_14633) );
CLKBUF_X2 inst_13194 ( .A(net_13041), .Z(net_13042) );
CLKBUF_X2 inst_10191 ( .A(net_10038), .Z(net_10039) );
AOI22_X2 inst_7794 ( .A2(net_6134), .B2(net_4809), .ZN(net_4795), .A1(net_4671), .B1(net_2501) );
CLKBUF_X2 inst_13349 ( .A(net_13196), .Z(net_13197) );
CLKBUF_X2 inst_17164 ( .A(net_14279), .Z(net_17012) );
CLKBUF_X2 inst_9355 ( .A(net_9202), .Z(net_9203) );
AOI221_X2 inst_8788 ( .ZN(net_5461), .B2(net_4973), .B1(net_853), .A(net_703), .C1(x12843), .C2(x1107) );
CLKBUF_X2 inst_16968 ( .A(net_16815), .Z(net_16816) );
CLKBUF_X2 inst_10128 ( .A(net_9491), .Z(net_9976) );
CLKBUF_X2 inst_10204 ( .A(net_10037), .Z(net_10052) );
NOR4_X2 inst_3217 ( .ZN(net_5735), .A1(net_5714), .A4(net_5712), .A2(net_5674), .A3(net_1532) );
CLKBUF_X2 inst_9556 ( .A(net_9403), .Z(net_9404) );
INV_X2 inst_6440 ( .ZN(net_627), .A(net_626) );
CLKBUF_X2 inst_14506 ( .A(net_14353), .Z(net_14354) );
NAND2_X2 inst_4376 ( .A1(net_7075), .A2(net_5162), .ZN(net_5081) );
CLKBUF_X2 inst_11778 ( .A(net_11625), .Z(net_11626) );
INV_X4 inst_6023 ( .A(net_5958), .ZN(x2633) );
CLKBUF_X2 inst_17845 ( .A(net_17692), .Z(net_17693) );
CLKBUF_X2 inst_18547 ( .A(net_10941), .Z(net_18395) );
OAI21_X2 inst_3044 ( .B2(net_8233), .B1(net_4928), .ZN(net_4778), .A(net_3206) );
INV_X4 inst_5443 ( .ZN(net_2669), .A(net_817) );
CLKBUF_X2 inst_14493 ( .A(net_13956), .Z(net_14341) );
CLKBUF_X2 inst_11914 ( .A(net_11761), .Z(net_11762) );
CLKBUF_X2 inst_12324 ( .A(net_12171), .Z(net_12172) );
SDFF_X2 inst_1072 ( .D(net_7311), .SI(net_6487), .Q(net_6487), .SE(net_3071), .CK(net_9929) );
SDFF_X2 inst_1993 ( .SI(net_7940), .Q(net_7940), .D(net_2656), .SE(net_2461), .CK(net_13992) );
CLKBUF_X2 inst_15744 ( .A(net_12498), .Z(net_15592) );
CLKBUF_X2 inst_14193 ( .A(net_14040), .Z(net_14041) );
CLKBUF_X2 inst_9791 ( .A(net_9638), .Z(net_9639) );
CLKBUF_X2 inst_15439 ( .A(net_15286), .Z(net_15287) );
HA_X1 inst_6671 ( .A(net_3332), .S(net_3199), .CO(net_3198), .B(net_3021) );
CLKBUF_X2 inst_17326 ( .A(net_17173), .Z(net_17174) );
CLKBUF_X2 inst_15580 ( .A(net_14021), .Z(net_15428) );
INV_X2 inst_6470 ( .A(net_7416), .ZN(net_572) );
NOR2_X2 inst_3617 ( .A1(net_5977), .A2(net_5976), .ZN(net_1101) );
CLKBUF_X2 inst_10893 ( .A(net_10740), .Z(net_10741) );
SDFF_X2 inst_1377 ( .SI(net_7274), .Q(net_7131), .D(net_7131), .SE(net_6279), .CK(net_14146) );
CLKBUF_X2 inst_15513 ( .A(net_15360), .Z(net_15361) );
CLKBUF_X2 inst_14828 ( .A(net_14141), .Z(net_14676) );
SDFFR_X2 inst_2201 ( .Q(net_7215), .D(net_2861), .SI(net_2843), .SE(net_1379), .CK(net_16141), .RN(x6501) );
CLKBUF_X2 inst_10581 ( .A(net_9080), .Z(net_10429) );
CLKBUF_X2 inst_14144 ( .A(net_13991), .Z(net_13992) );
CLKBUF_X2 inst_15835 ( .A(net_15682), .Z(net_15683) );
INV_X4 inst_5671 ( .A(net_8971), .ZN(net_1518) );
CLKBUF_X2 inst_17084 ( .A(net_12807), .Z(net_16932) );
CLKBUF_X2 inst_15990 ( .A(net_15837), .Z(net_15838) );
NAND2_X1 inst_4911 ( .A2(net_8268), .A1(net_6155), .ZN(net_730) );
NAND2_X2 inst_4525 ( .A1(net_3568), .ZN(net_3564), .A2(net_3563) );
NAND2_X2 inst_4115 ( .ZN(net_5413), .A1(net_5233), .A2(net_5009) );
CLKBUF_X2 inst_13264 ( .A(net_13111), .Z(net_13112) );
AOI22_X2 inst_8174 ( .B1(net_8789), .A1(net_8530), .ZN(net_6244), .A2(net_3861), .B2(net_3860) );
AOI22_X2 inst_8417 ( .B1(net_6718), .A1(net_6685), .B2(net_6202), .ZN(net_3525), .A2(net_3520) );
INV_X4 inst_5591 ( .A(net_6332), .ZN(net_689) );
SDFF_X2 inst_1687 ( .Q(net_8031), .D(net_8031), .SI(net_2713), .SE(net_2545), .CK(net_16470) );
CLKBUF_X2 inst_14983 ( .A(net_14830), .Z(net_14831) );
SDFF_X2 inst_1970 ( .D(net_7265), .SI(net_7002), .Q(net_7002), .SE(net_6277), .CK(net_17046) );
DFFR_X2 inst_7137 ( .QN(net_7352), .D(net_2987), .CK(net_9645), .RN(x6501) );
CLKBUF_X2 inst_12211 ( .A(net_12058), .Z(net_12059) );
DFF_X1 inst_6790 ( .Q(net_8251), .D(net_4428), .CK(net_16276) );
CLKBUF_X2 inst_14100 ( .A(net_13834), .Z(net_13948) );
CLKBUF_X2 inst_10256 ( .A(net_10103), .Z(net_10104) );
DFFR_X1 inst_7417 ( .D(net_5670), .CK(net_16763), .RN(x6501), .Q(x521) );
CLKBUF_X2 inst_12576 ( .A(net_12423), .Z(net_12424) );
NAND2_X2 inst_4842 ( .A1(net_8964), .A2(net_1887), .ZN(net_1103) );
SDFFR_X1 inst_2663 ( .D(net_6757), .SE(net_4506), .CK(net_9329), .RN(x6501), .SI(x2169), .Q(x2169) );
NOR3_X2 inst_3289 ( .A3(net_8953), .ZN(net_2237), .A1(net_2152), .A2(net_789) );
DFFR_X1 inst_7477 ( .QN(net_7429), .D(net_4220), .CK(net_12386), .RN(x6501) );
CLKBUF_X2 inst_15911 ( .A(net_15758), .Z(net_15759) );
CLKBUF_X2 inst_15597 ( .A(net_15444), .Z(net_15445) );
AOI22_X2 inst_7930 ( .B1(net_8180), .A1(net_7670), .B2(net_6099), .A2(net_4399), .ZN(net_4194) );
CLKBUF_X2 inst_12650 ( .A(net_12497), .Z(net_12498) );
CLKBUF_X2 inst_12116 ( .A(net_9416), .Z(net_11964) );
CLKBUF_X2 inst_10508 ( .A(net_10355), .Z(net_10356) );
CLKBUF_X2 inst_12087 ( .A(net_10605), .Z(net_11935) );
SDFF_X2 inst_401 ( .SI(net_8314), .Q(net_8314), .SE(net_3978), .D(net_3967), .CK(net_12291) );
AOI22_X2 inst_8086 ( .B1(net_8210), .A1(net_7700), .B2(net_6099), .A2(net_4399), .ZN(net_4060) );
OAI211_X2 inst_3210 ( .ZN(net_2118), .A(net_1894), .B(net_1853), .C1(net_1570), .C2(net_810) );
INV_X4 inst_5200 ( .A(net_5871), .ZN(net_5755) );
INV_X4 inst_6145 ( .A(net_6140), .ZN(net_6139) );
NAND2_X2 inst_4653 ( .ZN(net_2650), .A2(net_2649), .A1(net_1098) );
INV_X4 inst_6087 ( .A(net_7402), .ZN(net_701) );
CLKBUF_X2 inst_12028 ( .A(net_9217), .Z(net_11876) );
CLKBUF_X2 inst_17466 ( .A(net_9796), .Z(net_17314) );
CLKBUF_X2 inst_14823 ( .A(net_13430), .Z(net_14671) );
CLKBUF_X2 inst_18630 ( .A(net_18477), .Z(net_18478) );
NAND2_X2 inst_4465 ( .A2(net_4783), .ZN(net_4782), .A1(x1174) );
CLKBUF_X2 inst_13107 ( .A(net_9171), .Z(net_12955) );
CLKBUF_X2 inst_12281 ( .A(net_9232), .Z(net_12129) );
NAND2_X2 inst_4865 ( .A2(net_6169), .ZN(net_836), .A1(net_771) );
CLKBUF_X2 inst_13479 ( .A(net_13326), .Z(net_13327) );
AOI22_X2 inst_8548 ( .B1(net_6529), .A1(net_6496), .A2(net_6137), .B2(net_6104), .ZN(net_3392) );
SDFF_X2 inst_930 ( .SI(net_8717), .Q(net_8717), .SE(net_6195), .D(net_3966), .CK(net_12321) );
CLKBUF_X2 inst_11908 ( .A(net_9897), .Z(net_11756) );
DFF_X1 inst_6801 ( .QN(net_8220), .D(net_4432), .CK(net_17228) );
CLKBUF_X2 inst_15248 ( .A(net_15095), .Z(net_15096) );
AOI22_X2 inst_8494 ( .B1(net_6679), .A1(net_6646), .A2(net_6213), .B2(net_6138), .ZN(net_3446) );
CLKBUF_X2 inst_10453 ( .A(net_10300), .Z(net_10301) );
INV_X2 inst_6622 ( .A(net_6272), .ZN(net_6270) );
CLKBUF_X2 inst_18931 ( .A(net_18778), .Z(net_18779) );
CLKBUF_X2 inst_13650 ( .A(net_13497), .Z(net_13498) );
NAND3_X4 inst_3874 ( .A3(net_6057), .A1(net_6056), .ZN(net_2642), .A2(net_2094) );
AND2_X2 inst_9168 ( .A2(net_2554), .ZN(net_2552), .A1(net_2551) );
SDFF_X2 inst_1251 ( .SI(net_7696), .Q(net_7696), .SE(net_2714), .D(net_2710), .CK(net_13798) );
CLKBUF_X2 inst_12245 ( .A(net_10445), .Z(net_12093) );
DFFR_X2 inst_7360 ( .Q(net_7314), .CK(net_11373), .D(x13156), .RN(x6501) );
CLKBUF_X2 inst_12488 ( .A(net_11974), .Z(net_12336) );
CLKBUF_X2 inst_10300 ( .A(net_10147), .Z(net_10148) );
CLKBUF_X2 inst_10270 ( .A(net_10117), .Z(net_10118) );
DFFR_X1 inst_7433 ( .QN(net_8913), .D(net_4854), .CK(net_13984), .RN(x6501) );
CLKBUF_X2 inst_9937 ( .A(net_9784), .Z(net_9785) );
CLKBUF_X2 inst_18412 ( .A(net_9553), .Z(net_18260) );
CLKBUF_X2 inst_15411 ( .A(net_15112), .Z(net_15259) );
DFFR_X1 inst_7369 ( .D(net_5931), .CK(net_13912), .RN(x6501), .Q(x594) );
SDFFR_X2 inst_2172 ( .QN(net_7597), .SE(net_3144), .D(net_3129), .SI(net_1016), .CK(net_13506), .RN(x6501) );
AOI22_X2 inst_8005 ( .B1(net_7909), .A1(net_7807), .B2(net_6103), .A2(net_4398), .ZN(net_4129) );
SDFF_X2 inst_667 ( .Q(net_8442), .D(net_8442), .SI(net_3939), .SE(net_3934), .CK(net_12537) );
CLKBUF_X2 inst_15885 ( .A(net_15520), .Z(net_15733) );
CLKBUF_X2 inst_12646 ( .A(net_9843), .Z(net_12494) );
AOI21_X2 inst_8870 ( .B1(net_6342), .A(net_6341), .ZN(net_5941), .B2(net_5940) );
OR2_X2 inst_2896 ( .A1(net_7206), .A2(net_2255), .ZN(net_1723) );
CLKBUF_X2 inst_17477 ( .A(net_17324), .Z(net_17325) );
AOI221_X4 inst_8732 ( .B1(net_8848), .C1(net_8367), .C2(net_6265), .B2(net_6253), .ZN(net_4334), .A(net_4241) );
SDFFR_X1 inst_2691 ( .SI(net_7550), .SE(net_5043), .CK(net_12744), .RN(x6501), .Q(x3925), .D(x3925) );
CLKBUF_X2 inst_14401 ( .A(net_14003), .Z(net_14249) );
INV_X2 inst_6311 ( .ZN(net_3893), .A(net_3590) );
SDFF_X2 inst_1511 ( .SI(net_7872), .Q(net_7872), .D(net_2656), .SE(net_2558), .CK(net_14017) );
DFFR_X1 inst_7543 ( .D(net_916), .Q(net_392), .CK(net_16599), .RN(x6501) );
CLKBUF_X2 inst_10777 ( .A(net_10624), .Z(net_10625) );
CLKBUF_X2 inst_17839 ( .A(net_17686), .Z(net_17687) );
AOI21_X2 inst_8977 ( .B1(net_8214), .ZN(net_2189), .A(net_2188), .B2(net_2187) );
INV_X16 inst_6645 ( .ZN(net_3878), .A(net_3337) );
NAND2_X2 inst_4243 ( .A1(net_6904), .A2(net_5247), .ZN(net_5217) );
CLKBUF_X2 inst_18126 ( .A(net_17973), .Z(net_17974) );
CLKBUF_X2 inst_14344 ( .A(net_13431), .Z(net_14192) );
CLKBUF_X2 inst_13659 ( .A(net_12989), .Z(net_13507) );
SDFF_X2 inst_1504 ( .SI(net_7864), .Q(net_7864), .D(net_2717), .SE(net_2558), .CK(net_17012) );
CLKBUF_X2 inst_17730 ( .A(net_17577), .Z(net_17578) );
NOR2_X2 inst_3403 ( .A2(net_6158), .ZN(net_3929), .A1(net_3928) );
CLKBUF_X2 inst_18878 ( .A(net_18725), .Z(net_18726) );
INV_X4 inst_5830 ( .A(net_7515), .ZN(net_3332) );
CLKBUF_X2 inst_9802 ( .A(net_9649), .Z(net_9650) );
CLKBUF_X2 inst_19088 ( .A(net_18654), .Z(net_18936) );
CLKBUF_X2 inst_18961 ( .A(net_17680), .Z(net_18809) );
AOI211_X2 inst_9006 ( .C2(net_5595), .ZN(net_5474), .A(net_4948), .B(net_4936), .C1(net_323) );
DFFR_X1 inst_7518 ( .Q(net_302), .D(net_299), .CK(net_16610), .RN(x6501) );
DFFR_X2 inst_7242 ( .QN(net_7228), .D(net_2058), .CK(net_17788), .RN(x6501) );
NAND4_X2 inst_3807 ( .ZN(net_3619), .A1(net_3459), .A2(net_3458), .A3(net_3457), .A4(net_3456) );
CLKBUF_X2 inst_17825 ( .A(net_17672), .Z(net_17673) );
SDFF_X2 inst_1069 ( .D(net_7332), .SI(net_6541), .Q(net_6541), .SE(net_3086), .CK(net_9069) );
CLKBUF_X2 inst_12719 ( .A(net_12566), .Z(net_12567) );
CLKBUF_X2 inst_11327 ( .A(net_11174), .Z(net_11175) );
CLKBUF_X2 inst_18954 ( .A(net_18801), .Z(net_18802) );
CLKBUF_X2 inst_14153 ( .A(net_14000), .Z(net_14001) );
CLKBUF_X2 inst_13083 ( .A(net_12930), .Z(net_12931) );
CLKBUF_X2 inst_10326 ( .A(net_10173), .Z(net_10174) );
NOR2_X2 inst_3541 ( .ZN(net_1634), .A2(net_1481), .A1(net_1479) );
CLKBUF_X2 inst_11503 ( .A(net_11138), .Z(net_11351) );
CLKBUF_X2 inst_13825 ( .A(net_10287), .Z(net_13673) );
CLKBUF_X2 inst_17744 ( .A(net_17591), .Z(net_17592) );
INV_X4 inst_5167 ( .ZN(net_3294), .A(net_3031) );
NAND4_X2 inst_3850 ( .ZN(net_1620), .A2(net_1619), .A3(net_1618), .A4(net_1617), .A1(net_757) );
CLKBUF_X2 inst_16678 ( .A(net_16525), .Z(net_16526) );
CLKBUF_X2 inst_16533 ( .A(net_16380), .Z(net_16381) );
CLKBUF_X2 inst_12582 ( .A(net_9066), .Z(net_12430) );
CLKBUF_X2 inst_14368 ( .A(net_14215), .Z(net_14216) );
CLKBUF_X2 inst_10972 ( .A(net_10819), .Z(net_10820) );
SDFF_X2 inst_1786 ( .D(net_7301), .SI(net_6918), .Q(net_6918), .SE(net_6284), .CK(net_15885) );
CLKBUF_X2 inst_15271 ( .A(net_13366), .Z(net_15119) );
CLKBUF_X2 inst_15688 ( .A(net_15535), .Z(net_15536) );
SDFF_X2 inst_496 ( .SI(net_8622), .Q(net_8622), .SE(net_3984), .D(net_3952), .CK(net_10373) );
CLKBUF_X2 inst_10639 ( .A(net_10486), .Z(net_10487) );
DFFR_X2 inst_7174 ( .QN(net_7484), .D(net_2521), .CK(net_11214), .RN(x6501) );
CLKBUF_X2 inst_12356 ( .A(net_12203), .Z(net_12204) );
CLKBUF_X2 inst_10304 ( .A(net_10151), .Z(net_10152) );
INV_X4 inst_5369 ( .ZN(net_2796), .A(net_1361) );
CLKBUF_X2 inst_16889 ( .A(net_16736), .Z(net_16737) );
AOI211_X2 inst_9011 ( .C2(net_5267), .ZN(net_5047), .A(net_4905), .B(net_4734), .C1(net_166) );
INV_X4 inst_5733 ( .A(net_8929), .ZN(net_4518) );
DFFS_X2 inst_6867 ( .QN(net_7519), .D(net_4897), .CK(net_17619), .SN(x6501) );
NAND4_X2 inst_3749 ( .ZN(net_4281), .A1(net_4020), .A2(net_4019), .A3(net_4018), .A4(net_4017) );
SDFFR_X2 inst_2620 ( .Q(net_7371), .D(net_7371), .SE(net_1136), .CK(net_18621), .RN(x6501), .SI(x4812) );
CLKBUF_X2 inst_17115 ( .A(net_16962), .Z(net_16963) );
SDFF_X2 inst_1633 ( .Q(net_8178), .D(net_8178), .SI(net_2656), .SE(net_2538), .CK(net_14403) );
CLKBUF_X2 inst_12425 ( .A(net_11879), .Z(net_12273) );
SDFF_X2 inst_1262 ( .Q(net_8080), .D(net_8080), .SE(net_2707), .SI(net_2705), .CK(net_18580) );
INV_X4 inst_5303 ( .A(net_1662), .ZN(net_1621) );
CLKBUF_X2 inst_9364 ( .A(net_9168), .Z(net_9212) );
AOI22_X2 inst_8048 ( .B1(net_8035), .A1(net_8001), .B2(net_6102), .A2(net_6097), .ZN(net_4092) );
CLKBUF_X2 inst_16882 ( .A(net_16729), .Z(net_16730) );
DFF_X1 inst_6799 ( .Q(net_8246), .D(net_4434), .CK(net_16273) );
NAND4_X2 inst_3856 ( .A1(net_6382), .A4(net_6380), .A3(net_1492), .ZN(net_1259), .A2(net_1258) );
CLKBUF_X2 inst_12453 ( .A(net_12300), .Z(net_12301) );
INV_X4 inst_5091 ( .ZN(net_5706), .A(net_5682) );
CLKBUF_X2 inst_14169 ( .A(net_14016), .Z(net_14017) );
CLKBUF_X2 inst_11650 ( .A(net_10343), .Z(net_11498) );
CLKBUF_X2 inst_12577 ( .A(net_12253), .Z(net_12425) );
CLKBUF_X2 inst_11482 ( .A(net_10242), .Z(net_11330) );
INV_X2 inst_6432 ( .ZN(net_696), .A(net_695) );
CLKBUF_X2 inst_16891 ( .A(net_16738), .Z(net_16739) );
CLKBUF_X2 inst_10716 ( .A(net_10563), .Z(net_10564) );
CLKBUF_X2 inst_16615 ( .A(net_14480), .Z(net_16463) );
SDFF_X2 inst_1077 ( .D(net_7327), .SI(net_6503), .Q(net_6503), .SE(net_3071), .CK(net_9854) );
CLKBUF_X2 inst_15495 ( .A(net_14962), .Z(net_15343) );
INV_X2 inst_6461 ( .A(net_6473), .ZN(net_3284) );
SDFFR_X1 inst_2757 ( .QN(net_7589), .D(net_3953), .SE(net_3144), .SI(net_623), .CK(net_12573), .RN(x6501) );
SDFF_X2 inst_1932 ( .SI(net_8062), .Q(net_8062), .D(net_2590), .SE(net_2508), .CK(net_15954) );
CLKBUF_X2 inst_10822 ( .A(net_10532), .Z(net_10670) );
CLKBUF_X2 inst_9733 ( .A(net_9580), .Z(net_9581) );
AOI22_X2 inst_7884 ( .A2(net_5538), .ZN(net_4547), .B2(net_4388), .B1(net_2596), .A1(net_424) );
NAND4_X2 inst_3704 ( .ZN(net_4433), .A4(net_4337), .A1(net_3740), .A2(net_3739), .A3(net_3738) );
CLKBUF_X2 inst_13903 ( .A(net_13750), .Z(net_13751) );
CLKBUF_X2 inst_11828 ( .A(net_11675), .Z(net_11676) );
CLKBUF_X2 inst_18792 ( .A(net_18639), .Z(net_18640) );
CLKBUF_X2 inst_17129 ( .A(net_16976), .Z(net_16977) );
SDFF_X2 inst_1052 ( .SI(net_7332), .Q(net_6673), .D(net_6673), .SE(net_3126), .CK(net_9073) );
SDFF_X2 inst_1280 ( .Q(net_8082), .D(net_8082), .SI(net_2709), .SE(net_2707), .CK(net_15780) );
CLKBUF_X2 inst_12740 ( .A(net_9058), .Z(net_12588) );
INV_X2 inst_6435 ( .ZN(net_684), .A(net_683) );
INV_X4 inst_5362 ( .ZN(net_1141), .A(net_1140) );
CLKBUF_X2 inst_13904 ( .A(net_13751), .Z(net_13752) );
CLKBUF_X2 inst_9578 ( .A(net_9425), .Z(net_9426) );
INV_X4 inst_6112 ( .A(net_6409), .ZN(net_1843) );
INV_X2 inst_6200 ( .ZN(net_5510), .A(net_5429) );
CLKBUF_X2 inst_14975 ( .A(net_10437), .Z(net_14823) );
CLKBUF_X2 inst_16513 ( .A(net_16360), .Z(net_16361) );
XNOR2_X2 inst_134 ( .B(net_7616), .ZN(net_2812), .A(net_2497) );
SDFFR_X2 inst_2409 ( .SI(net_5945), .SE(net_2260), .Q(net_348), .D(net_348), .CK(net_9352), .RN(x6501) );
NOR2_X4 inst_3322 ( .ZN(net_6254), .A1(net_5591), .A2(net_5589) );
NOR2_X2 inst_3425 ( .ZN(net_3092), .A1(net_3023), .A2(net_2984) );
SDFFR_X2 inst_2328 ( .SI(net_7366), .D(net_2742), .SE(net_2740), .QN(net_277), .CK(net_13696), .RN(x6501) );
AOI22_X2 inst_8060 ( .B1(net_8071), .A1(net_7867), .B2(net_6107), .A2(net_4400), .ZN(net_4082) );
INV_X4 inst_5779 ( .A(net_7193), .ZN(net_2955) );
CLKBUF_X2 inst_14890 ( .A(net_14737), .Z(net_14738) );
CLKBUF_X2 inst_18285 ( .A(net_18132), .Z(net_18133) );
CLKBUF_X2 inst_13541 ( .A(net_13388), .Z(net_13389) );
OAI22_X2 inst_2912 ( .A1(net_4922), .ZN(net_4775), .B2(net_4774), .A2(net_4511), .B1(net_1799) );
SDFF_X2 inst_762 ( .Q(net_8804), .D(net_8804), .SI(net_3975), .SE(net_3879), .CK(net_12521) );
OAI21_X2 inst_3025 ( .B2(net_4971), .ZN(net_4967), .A(net_4804), .B1(net_624) );
CLKBUF_X2 inst_15472 ( .A(net_15319), .Z(net_15320) );
CLKBUF_X2 inst_15600 ( .A(net_15447), .Z(net_15448) );
DFFR_X1 inst_7530 ( .Q(net_6468), .D(net_6465), .CK(net_15131), .RN(x6501) );
CLKBUF_X2 inst_16649 ( .A(net_16496), .Z(net_16497) );
CLKBUF_X2 inst_10434 ( .A(net_10281), .Z(net_10282) );
CLKBUF_X2 inst_16171 ( .A(net_16018), .Z(net_16019) );
NAND2_X2 inst_4530 ( .ZN(net_3383), .A2(net_3381), .A1(net_3367) );
CLKBUF_X2 inst_11882 ( .A(net_10327), .Z(net_11730) );
CLKBUF_X2 inst_14607 ( .A(net_10490), .Z(net_14455) );
CLKBUF_X2 inst_13843 ( .A(net_13690), .Z(net_13691) );
SDFF_X2 inst_1956 ( .D(net_7289), .SI(net_7026), .Q(net_7026), .SE(net_6277), .CK(net_18357) );
AOI22_X2 inst_8378 ( .B1(net_8782), .A1(net_8523), .A2(net_3861), .B2(net_3860), .ZN(net_3670) );
CLKBUF_X2 inst_10687 ( .A(net_10534), .Z(net_10535) );
CLKBUF_X2 inst_10935 ( .A(net_10782), .Z(net_10783) );
SDFF_X2 inst_751 ( .Q(net_8791), .D(net_8791), .SI(net_3966), .SE(net_3879), .CK(net_10905) );
CLKBUF_X2 inst_19195 ( .A(net_19042), .Z(net_19043) );
NAND2_X2 inst_4283 ( .A1(net_6886), .A2(net_5247), .ZN(net_5177) );
SDFFR_X2 inst_2471 ( .SE(net_2678), .D(net_2570), .SI(net_436), .Q(net_436), .CK(net_14811), .RN(x6501) );
NOR4_X2 inst_3244 ( .ZN(net_1559), .A1(net_1094), .A2(net_993), .A3(net_952), .A4(net_950) );
NAND4_X2 inst_3821 ( .ZN(net_3605), .A1(net_3403), .A2(net_3402), .A3(net_3401), .A4(net_3400) );
DFFR_X1 inst_7443 ( .QN(net_8923), .D(net_4760), .CK(net_17317), .RN(x6501) );
INV_X4 inst_5981 ( .A(net_6356), .ZN(net_513) );
CLKBUF_X2 inst_14554 ( .A(net_12647), .Z(net_14402) );
CLKBUF_X2 inst_12675 ( .A(net_12522), .Z(net_12523) );
CLKBUF_X2 inst_13330 ( .A(net_9570), .Z(net_13178) );
NAND2_X2 inst_4623 ( .A2(net_6144), .ZN(net_2595), .A1(net_2594) );
NAND4_X2 inst_3835 ( .ZN(net_2111), .A4(net_1831), .A3(net_1647), .A1(net_1040), .A2(net_995) );
SDFFR_X2 inst_2117 ( .SI(net_7200), .Q(net_7200), .D(net_6451), .SE(net_4362), .CK(net_14570), .RN(x6501) );
OAI21_X2 inst_3140 ( .B1(net_5957), .B2(net_2060), .ZN(net_2057), .A(net_2056) );
CLKBUF_X2 inst_13812 ( .A(net_13659), .Z(net_13660) );
CLKBUF_X2 inst_12035 ( .A(net_11882), .Z(net_11883) );
CLKBUF_X2 inst_17775 ( .A(net_12144), .Z(net_17623) );
CLKBUF_X2 inst_14600 ( .A(net_9154), .Z(net_14448) );
CLKBUF_X2 inst_11941 ( .A(net_9878), .Z(net_11789) );
CLKBUF_X2 inst_12308 ( .A(net_11584), .Z(net_12156) );
CLKBUF_X2 inst_11200 ( .A(net_9190), .Z(net_11048) );
NAND2_X2 inst_4642 ( .ZN(net_2801), .A2(net_2418), .A1(net_2113) );
DFFR_X2 inst_7340 ( .Q(net_7317), .CK(net_11385), .D(x13126), .RN(x6501) );
NOR3_X2 inst_3316 ( .A2(net_7399), .ZN(net_4275), .A1(net_1369), .A3(net_867) );
CLKBUF_X2 inst_19051 ( .A(net_17690), .Z(net_18899) );
CLKBUF_X2 inst_9385 ( .A(net_9100), .Z(net_9233) );
NAND2_X2 inst_4411 ( .A1(net_6850), .ZN(net_5017), .A2(net_5016) );
CLKBUF_X2 inst_11471 ( .A(net_11318), .Z(net_11319) );
AOI22_X2 inst_7772 ( .B1(net_6999), .A1(net_6959), .A2(net_5443), .B2(net_5442), .ZN(net_5315) );
NAND2_X4 inst_4014 ( .ZN(net_4456), .A1(net_4375), .A2(net_4361) );
CLKBUF_X2 inst_17087 ( .A(net_14425), .Z(net_16935) );
NAND4_X2 inst_3694 ( .ZN(net_4443), .A4(net_4343), .A1(net_3800), .A2(net_3799), .A3(net_3798) );
CLKBUF_X2 inst_16272 ( .A(net_16119), .Z(net_16120) );
CLKBUF_X2 inst_15204 ( .A(net_12075), .Z(net_15052) );
NAND2_X2 inst_4882 ( .A2(net_7393), .ZN(net_775), .A1(net_182) );
SDFFR_X1 inst_2698 ( .SI(net_7530), .SE(net_5043), .CK(net_11946), .RN(x6501), .Q(x4179), .D(x4179) );
CLKBUF_X2 inst_9908 ( .A(net_9244), .Z(net_9756) );
SDFFR_X2 inst_2518 ( .D(net_7378), .SE(net_2376), .SI(net_211), .Q(net_211), .CK(net_17751), .RN(x6501) );
NOR2_X2 inst_3460 ( .A2(net_3080), .ZN(net_2782), .A1(net_2781) );
INV_X4 inst_5152 ( .ZN(net_3259), .A(net_3221) );
INV_X4 inst_5544 ( .ZN(net_826), .A(net_644) );
SDFFS_X2 inst_2075 ( .SI(net_7375), .SE(net_2794), .Q(net_164), .D(net_164), .CK(net_17736), .SN(x6501) );
SDFF_X2 inst_1911 ( .D(net_7278), .SI(net_6895), .Q(net_6895), .SE(net_6284), .CK(net_14601) );
INV_X4 inst_5689 ( .ZN(net_2695), .A(net_147) );
CLKBUF_X2 inst_10841 ( .A(net_10065), .Z(net_10689) );
CLKBUF_X2 inst_15528 ( .A(net_12167), .Z(net_15376) );
SDFF_X2 inst_585 ( .Q(net_8819), .D(net_8819), .SE(net_3964), .SI(net_3938), .CK(net_10733) );
CLKBUF_X2 inst_15846 ( .A(net_12126), .Z(net_15694) );
AOI221_X2 inst_8816 ( .C2(net_5535), .B2(net_5260), .A(net_4898), .ZN(net_4711), .B1(net_3205), .C1(net_459) );
INV_X4 inst_5435 ( .ZN(net_1142), .A(net_826) );
INV_X4 inst_5107 ( .ZN(net_4953), .A(net_4900) );
INV_X4 inst_5763 ( .A(net_7593), .ZN(net_2836) );
CLKBUF_X2 inst_11171 ( .A(net_10384), .Z(net_11019) );
CLKBUF_X2 inst_18428 ( .A(net_9692), .Z(net_18276) );
CLKBUF_X2 inst_12137 ( .A(net_11984), .Z(net_11985) );
INV_X2 inst_6453 ( .A(net_6476), .ZN(net_589) );
SDFFR_X2 inst_2428 ( .SE(net_2683), .D(net_2673), .SI(net_451), .Q(net_451), .CK(net_13841), .RN(x6501) );
INV_X4 inst_5115 ( .ZN(net_4783), .A(net_4642) );
CLKBUF_X2 inst_14382 ( .A(net_12854), .Z(net_14230) );
DFFR_X1 inst_7553 ( .D(net_2697), .Q(net_292), .CK(net_11629), .RN(x6501) );
CLKBUF_X2 inst_18966 ( .A(net_18813), .Z(net_18814) );
CLKBUF_X2 inst_17264 ( .A(net_9408), .Z(net_17112) );
SDFF_X2 inst_1124 ( .D(net_7330), .SI(net_6572), .Q(net_6572), .SE(net_3070), .CK(net_11311) );
NAND2_X2 inst_4086 ( .ZN(net_5747), .A1(net_5691), .A2(net_5688) );
CLKBUF_X2 inst_11091 ( .A(net_9186), .Z(net_10939) );
SDFFR_X2 inst_2555 ( .QN(net_6378), .SE(net_2147), .SI(net_1939), .D(net_948), .CK(net_15355), .RN(x6501) );
CLKBUF_X2 inst_13922 ( .A(net_13769), .Z(net_13770) );
DFFS_X1 inst_6966 ( .D(net_6828), .Q(net_6801), .CK(net_9628), .SN(x6501) );
CLKBUF_X2 inst_18526 ( .A(net_9640), .Z(net_18374) );
CLKBUF_X2 inst_13447 ( .A(net_13294), .Z(net_13295) );
INV_X4 inst_5240 ( .ZN(net_2328), .A(net_2172) );
CLKBUF_X2 inst_12450 ( .A(net_12297), .Z(net_12298) );
INV_X4 inst_5343 ( .A(net_1836), .ZN(net_1288) );
NAND4_X2 inst_3714 ( .ZN(net_4423), .A4(net_4330), .A1(net_3673), .A2(net_3672), .A3(net_3671) );
CLKBUF_X2 inst_12317 ( .A(net_11468), .Z(net_12165) );
CLKBUF_X2 inst_12269 ( .A(net_12116), .Z(net_12117) );
INV_X4 inst_5285 ( .ZN(net_2048), .A(net_1379) );
CLKBUF_X2 inst_17972 ( .A(net_13716), .Z(net_17820) );
INV_X1 inst_6658 ( .A(net_6193), .ZN(net_6192) );
INV_X4 inst_5611 ( .A(net_6365), .ZN(net_697) );
SDFF_X2 inst_1304 ( .Q(net_7821), .D(net_7821), .SE(net_2730), .SI(net_2576), .CK(net_18889) );
AND4_X4 inst_9027 ( .A3(net_3227), .ZN(net_3192), .A2(net_3087), .A1(net_1441), .A4(net_537) );
DFF_X1 inst_6815 ( .QN(net_8230), .D(net_4451), .CK(net_17218) );
NOR3_X2 inst_3292 ( .A1(net_2400), .ZN(net_2339), .A3(net_2180), .A2(net_1876) );
AOI22_X2 inst_8575 ( .A2(net_1996), .ZN(net_1815), .A1(net_1814), .B1(net_1813), .B2(net_1812) );
AOI22_X2 inst_7751 ( .B1(net_6961), .A1(net_6921), .A2(net_5443), .B2(net_5442), .ZN(net_5402) );
INV_X8 inst_5024 ( .ZN(net_3978), .A(net_3329) );
SDFF_X2 inst_919 ( .SI(net_8740), .Q(net_8740), .SE(net_6195), .D(net_3948), .CK(net_13387) );
CLKBUF_X2 inst_10530 ( .A(net_10377), .Z(net_10378) );
CLKBUF_X2 inst_12772 ( .A(net_12619), .Z(net_12620) );
SDFF_X2 inst_1916 ( .D(net_7272), .SI(net_6929), .Q(net_6929), .SE(net_6281), .CK(net_14082) );
CLKBUF_X2 inst_9705 ( .A(net_9552), .Z(net_9553) );
CLKBUF_X2 inst_14057 ( .A(net_9596), .Z(net_13905) );
CLKBUF_X2 inst_12403 ( .A(net_11555), .Z(net_12251) );
SDFF_X2 inst_1797 ( .SI(net_8064), .Q(net_8064), .D(net_2718), .SE(net_2508), .CK(net_18758) );
CLKBUF_X2 inst_17447 ( .A(net_17294), .Z(net_17295) );
NAND2_X2 inst_4408 ( .A1(net_7089), .A2(net_5164), .ZN(net_5049) );
SDFFR_X1 inst_2708 ( .SI(net_6812), .Q(net_6812), .SE(net_6270), .D(net_6142), .CK(net_9619), .RN(x6501) );
INV_X2 inst_6197 ( .ZN(net_5513), .A(net_5441) );
CLKBUF_X2 inst_14694 ( .A(net_10936), .Z(net_14542) );
CLKBUF_X2 inst_9866 ( .A(net_9713), .Z(net_9714) );
NOR2_X2 inst_3530 ( .ZN(net_1683), .A2(net_1327), .A1(net_1138) );
INV_X8 inst_5009 ( .ZN(net_5535), .A(net_4470) );
NAND2_X2 inst_4785 ( .A1(net_2207), .ZN(net_1730), .A2(net_1535) );
CLKBUF_X2 inst_13552 ( .A(net_12245), .Z(net_13400) );
AOI22_X2 inst_7785 ( .A1(net_5268), .ZN(net_4865), .B2(net_4809), .A2(net_4630), .B1(net_350) );
SDFFR_X2 inst_2592 ( .D(net_7390), .QN(net_7250), .SI(net_1944), .SE(net_1379), .CK(net_18107), .RN(x6501) );
CLKBUF_X2 inst_18297 ( .A(net_18144), .Z(net_18145) );
CLKBUF_X2 inst_12752 ( .A(net_12599), .Z(net_12600) );
DFFR_X2 inst_7331 ( .D(net_7171), .QN(net_7169), .CK(net_9557), .RN(x6501) );
OAI21_X2 inst_3116 ( .A(net_2473), .ZN(net_2410), .B2(net_2327), .B1(net_2171) );
CLKBUF_X2 inst_17106 ( .A(net_16953), .Z(net_16954) );
CLKBUF_X2 inst_15624 ( .A(net_15471), .Z(net_15472) );
NAND2_X2 inst_4378 ( .A1(net_7116), .A2(net_5164), .ZN(net_5079) );
CLKBUF_X2 inst_14682 ( .A(net_14529), .Z(net_14530) );
CLKBUF_X2 inst_9682 ( .A(net_9067), .Z(net_9530) );
CLKBUF_X2 inst_15824 ( .A(net_15671), .Z(net_15672) );
CLKBUF_X2 inst_15589 ( .A(net_15436), .Z(net_15437) );
CLKBUF_X2 inst_15552 ( .A(net_15399), .Z(net_15400) );
XNOR2_X2 inst_114 ( .ZN(net_3547), .B(net_3546), .A(net_3276) );
CLKBUF_X2 inst_11767 ( .A(net_10198), .Z(net_11615) );
DFFR_X2 inst_7116 ( .QN(net_7613), .D(net_3054), .CK(net_9807), .RN(x6501) );
SDFFR_X2 inst_2278 ( .SI(net_2796), .SE(net_2789), .Q(net_250), .D(net_250), .CK(net_18333), .RN(x6501) );
NAND2_X2 inst_4866 ( .A1(net_7165), .ZN(net_1922), .A2(net_835) );
CLKBUF_X2 inst_11415 ( .A(net_11262), .Z(net_11263) );
AOI22_X2 inst_7924 ( .B1(net_8146), .A1(net_7704), .B2(net_6101), .A2(net_6095), .ZN(net_5996) );
AOI22_X2 inst_7800 ( .A2(net_6130), .B2(net_4965), .ZN(net_4788), .A1(net_1425), .B1(net_306) );
NAND2_X2 inst_4150 ( .ZN(net_5367), .A2(net_5210), .A1(net_5105) );
CLKBUF_X2 inst_9630 ( .A(net_9420), .Z(net_9478) );
CLKBUF_X2 inst_12371 ( .A(net_12218), .Z(net_12219) );
SDFF_X2 inst_534 ( .Q(net_8859), .D(net_8859), .SI(net_3981), .SE(net_3936), .CK(net_12454) );
CLKBUF_X2 inst_12422 ( .A(net_12269), .Z(net_12270) );
CLKBUF_X2 inst_16879 ( .A(net_9561), .Z(net_16727) );
AOI222_X1 inst_8636 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_4225), .B1(net_3534), .C1(net_3533), .A1(x13674) );
CLKBUF_X2 inst_17268 ( .A(net_17115), .Z(net_17116) );
CLKBUF_X2 inst_13816 ( .A(net_13663), .Z(net_13664) );
CLKBUF_X2 inst_18679 ( .A(net_18526), .Z(net_18527) );
AND4_X2 inst_9033 ( .ZN(net_5606), .A2(net_5536), .A1(net_4868), .A3(net_4544), .A4(net_4543) );
CLKBUF_X2 inst_16476 ( .A(net_16323), .Z(net_16324) );
CLKBUF_X2 inst_10682 ( .A(net_10529), .Z(net_10530) );
INV_X4 inst_5618 ( .A(net_8922), .ZN(net_2626) );
CLKBUF_X2 inst_18632 ( .A(net_17062), .Z(net_18480) );
CLKBUF_X2 inst_15318 ( .A(net_15165), .Z(net_15166) );
INV_X4 inst_5193 ( .ZN(net_2847), .A(net_2799) );
OR2_X4 inst_2836 ( .ZN(net_6144), .A2(net_2482), .A1(net_1724) );
NAND2_X2 inst_4336 ( .A1(net_7103), .A2(net_5164), .ZN(net_5121) );
CLKBUF_X2 inst_17350 ( .A(net_14730), .Z(net_17198) );
CLKBUF_X2 inst_16448 ( .A(net_15424), .Z(net_16296) );
CLKBUF_X2 inst_18227 ( .A(net_18074), .Z(net_18075) );
CLKBUF_X2 inst_10424 ( .A(net_10271), .Z(net_10272) );
SDFFR_X1 inst_2770 ( .D(net_7390), .Q(net_7287), .SI(net_1944), .SE(net_1327), .CK(net_18171), .RN(x6501) );
CLKBUF_X2 inst_11735 ( .A(net_11582), .Z(net_11583) );
AND2_X2 inst_9184 ( .ZN(net_2140), .A1(net_1949), .A2(net_1948) );
CLKBUF_X2 inst_14542 ( .A(net_14389), .Z(net_14390) );
CLKBUF_X2 inst_15010 ( .A(net_14857), .Z(net_14858) );
NAND2_X2 inst_4573 ( .ZN(net_2998), .A1(net_2997), .A2(net_2996) );
NOR2_X2 inst_3444 ( .A2(net_3093), .ZN(net_3044), .A1(net_2227) );
DFFR_X2 inst_7284 ( .Q(net_9008), .D(net_1726), .CK(net_16288), .RN(x6501) );
CLKBUF_X2 inst_10848 ( .A(net_9831), .Z(net_10696) );
CLKBUF_X2 inst_9295 ( .A(net_9142), .Z(net_9143) );
CLKBUF_X2 inst_14926 ( .A(net_14773), .Z(net_14774) );
NAND2_X2 inst_4732 ( .ZN(net_2573), .A2(net_1586), .A1(net_930) );
CLKBUF_X2 inst_17655 ( .A(net_13104), .Z(net_17503) );
SDFFR_X2 inst_2348 ( .SI(net_7367), .D(net_2733), .SE(net_2732), .QN(net_271), .CK(net_16128), .RN(x6501) );
NAND2_X4 inst_4021 ( .A1(net_6158), .ZN(net_4216), .A2(net_2847) );
CLKBUF_X2 inst_11059 ( .A(net_10906), .Z(net_10907) );
CLKBUF_X2 inst_9827 ( .A(net_9674), .Z(net_9675) );
CLKBUF_X2 inst_18421 ( .A(net_17146), .Z(net_18269) );
AOI22_X2 inst_8290 ( .A1(net_8619), .B1(net_8434), .A2(net_3864), .B2(net_3863), .ZN(net_3752) );
CLKBUF_X2 inst_11114 ( .A(net_10961), .Z(net_10962) );
INV_X4 inst_5080 ( .ZN(net_5760), .A(net_5724) );
NAND2_X2 inst_4666 ( .A2(net_2328), .ZN(net_2169), .A1(net_1663) );
CLKBUF_X2 inst_16104 ( .A(net_15951), .Z(net_15952) );
CLKBUF_X2 inst_14115 ( .A(net_13962), .Z(net_13963) );
SDFF_X2 inst_1465 ( .SI(net_7290), .Q(net_7147), .D(net_7147), .SE(net_6279), .CK(net_18278) );
INV_X4 inst_5265 ( .ZN(net_2129), .A(net_1932) );
CLKBUF_X2 inst_13009 ( .A(net_12856), .Z(net_12857) );
INV_X2 inst_6550 ( .A(net_6367), .ZN(net_2134) );
CLKBUF_X2 inst_17205 ( .A(net_17052), .Z(net_17053) );
CLKBUF_X2 inst_15069 ( .A(net_14916), .Z(net_14917) );
CLKBUF_X2 inst_18334 ( .A(net_18181), .Z(net_18182) );
NAND2_X2 inst_4215 ( .A1(net_6891), .A2(net_5247), .ZN(net_5245) );
CLKBUF_X2 inst_15259 ( .A(net_15106), .Z(net_15107) );
SDFF_X2 inst_999 ( .D(net_7339), .SI(net_6647), .Q(net_6647), .SE(net_3123), .CK(net_11910) );
AOI22_X2 inst_7805 ( .A2(net_8223), .B1(net_7179), .B2(net_5655), .A1(net_5268), .ZN(net_4769) );
CLKBUF_X2 inst_12378 ( .A(net_11713), .Z(net_12226) );
CLKBUF_X2 inst_19105 ( .A(net_15276), .Z(net_18953) );
AOI22_X2 inst_8083 ( .B1(net_8148), .A1(net_7706), .B2(net_6101), .A2(net_6095), .ZN(net_4062) );
SDFF_X2 inst_1846 ( .SI(net_6916), .Q(net_6916), .SE(net_6284), .D(net_2544), .CK(net_18666) );
SDFFR_X2 inst_2139 ( .SI(net_7198), .Q(net_7198), .D(net_6449), .SE(net_4362), .CK(net_16433), .RN(x6501) );
CLKBUF_X2 inst_17565 ( .A(net_17412), .Z(net_17413) );
NAND2_X2 inst_4278 ( .A1(net_7004), .A2(net_5249), .ZN(net_5182) );
CLKBUF_X2 inst_10236 ( .A(net_10083), .Z(net_10084) );
XNOR2_X2 inst_186 ( .A(net_7661), .ZN(net_1644), .B(net_1643) );
NAND2_X2 inst_4271 ( .A1(net_6917), .A2(net_5247), .ZN(net_5189) );
CLKBUF_X2 inst_16066 ( .A(net_12264), .Z(net_15914) );
CLKBUF_X2 inst_10756 ( .A(net_10603), .Z(net_10604) );
CLKBUF_X2 inst_9820 ( .A(net_9346), .Z(net_9668) );
OAI21_X2 inst_3071 ( .ZN(net_4226), .A(net_3883), .B2(net_3552), .B1(net_1375) );
CLKBUF_X2 inst_10395 ( .A(net_10242), .Z(net_10243) );
CLKBUF_X2 inst_11963 ( .A(net_11810), .Z(net_11811) );
CLKBUF_X2 inst_13536 ( .A(net_13383), .Z(net_13384) );
AOI22_X2 inst_8283 ( .B1(net_8877), .A1(net_8322), .B2(net_6252), .A2(net_4345), .ZN(net_3758) );
SDFF_X2 inst_863 ( .Q(net_8572), .D(net_8572), .SI(net_3944), .SE(net_3878), .CK(net_12246) );
CLKBUF_X2 inst_16821 ( .A(net_16668), .Z(net_16669) );
AOI222_X1 inst_8669 ( .A1(net_7649), .A2(net_3599), .B2(net_3598), .C2(net_3597), .ZN(net_3589), .C1(net_1643), .B1(net_526) );
INV_X2 inst_6315 ( .ZN(net_3348), .A(net_3297) );
SDFF_X2 inst_1385 ( .SI(net_7733), .Q(net_7733), .D(net_2660), .SE(net_2559), .CK(net_17015) );
CLKBUF_X2 inst_15288 ( .A(net_15135), .Z(net_15136) );
INV_X2 inst_6513 ( .A(net_8268), .ZN(net_533) );
INV_X4 inst_5921 ( .A(net_7247), .ZN(net_1957) );
INV_X4 inst_5770 ( .A(net_7226), .ZN(net_1615) );
SDFF_X2 inst_1573 ( .Q(net_8021), .D(net_8021), .SI(net_2706), .SE(net_2545), .CK(net_15271) );
INV_X4 inst_5521 ( .ZN(net_863), .A(net_672) );
AOI22_X2 inst_8394 ( .B1(net_8821), .A1(net_8340), .A2(net_6265), .B2(net_6253), .ZN(net_6070) );
SDFF_X2 inst_1390 ( .SI(net_7287), .Q(net_7104), .D(net_7104), .SE(net_6278), .CK(net_14930) );
CLKBUF_X2 inst_18738 ( .A(net_18585), .Z(net_18586) );
XNOR2_X2 inst_229 ( .ZN(net_1313), .A(net_1101), .B(net_885) );
AND2_X4 inst_9124 ( .A2(net_7405), .ZN(net_1376), .A1(net_717) );
CLKBUF_X2 inst_19008 ( .A(net_18855), .Z(net_18856) );
CLKBUF_X2 inst_12920 ( .A(net_12363), .Z(net_12768) );
CLKBUF_X2 inst_9596 ( .A(net_9215), .Z(net_9444) );
MUX2_X2 inst_4992 ( .A(net_9024), .Z(net_3946), .B(net_2462), .S(net_622) );
NAND2_X2 inst_4689 ( .ZN(net_6217), .A2(net_6157), .A1(net_808) );
CLKBUF_X2 inst_17063 ( .A(net_16910), .Z(net_16911) );
CLKBUF_X2 inst_11719 ( .A(net_9511), .Z(net_11567) );
INV_X4 inst_6151 ( .A(net_6179), .ZN(net_6178) );
AND2_X2 inst_9187 ( .A2(net_7620), .ZN(net_1842), .A1(net_1563) );
SDFFR_X2 inst_2131 ( .SI(net_7196), .Q(net_7196), .D(net_6447), .SE(net_4362), .CK(net_13560), .RN(x6501) );
CLKBUF_X2 inst_12007 ( .A(net_11854), .Z(net_11855) );
CLKBUF_X2 inst_9949 ( .A(net_9796), .Z(net_9797) );
DFFR_X2 inst_7297 ( .QN(net_7220), .D(net_1631), .CK(net_15179), .RN(x6501) );
AOI221_X2 inst_8804 ( .C2(net_8218), .B2(net_5520), .C1(net_5268), .A(net_4905), .ZN(net_4826), .B1(net_281) );
CLKBUF_X2 inst_9453 ( .A(net_9107), .Z(net_9301) );
SDFF_X2 inst_421 ( .SI(net_8303), .Q(net_8303), .SE(net_3978), .D(net_3947), .CK(net_13004) );
CLKBUF_X2 inst_11263 ( .A(net_10447), .Z(net_11111) );
DFFR_X2 inst_7016 ( .QN(net_6288), .D(net_5730), .CK(net_13878), .RN(x6501) );
SDFF_X2 inst_816 ( .SI(net_8507), .Q(net_8507), .D(net_3954), .SE(net_3884), .CK(net_10981) );
CLKBUF_X2 inst_11000 ( .A(net_10112), .Z(net_10848) );
CLKBUF_X2 inst_16824 ( .A(net_16671), .Z(net_16672) );
CLKBUF_X2 inst_12911 ( .A(net_12608), .Z(net_12759) );
OR3_X4 inst_2798 ( .A2(net_6126), .ZN(net_2952), .A3(net_2526), .A1(net_2348) );
CLKBUF_X2 inst_12903 ( .A(net_12750), .Z(net_12751) );
CLKBUF_X2 inst_12692 ( .A(net_10796), .Z(net_12540) );
CLKBUF_X2 inst_13694 ( .A(net_13541), .Z(net_13542) );
SDFF_X2 inst_1108 ( .D(net_7339), .SI(net_6548), .Q(net_6548), .SE(net_3086), .CK(net_11874) );
CLKBUF_X2 inst_19013 ( .A(net_18860), .Z(net_18861) );
INV_X4 inst_5148 ( .A(net_3887), .ZN(net_3597) );
NAND2_X2 inst_4534 ( .A1(net_3381), .ZN(net_3377), .A2(net_3369) );
AOI22_X2 inst_8286 ( .B1(net_8804), .A1(net_8545), .A2(net_3861), .B2(net_3860), .ZN(net_3756) );
CLKBUF_X2 inst_15901 ( .A(net_15748), .Z(net_15749) );
CLKBUF_X2 inst_11422 ( .A(net_11269), .Z(net_11270) );
CLKBUF_X2 inst_16288 ( .A(net_16135), .Z(net_16136) );
AOI222_X1 inst_8604 ( .B2(net_6770), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5820), .A1(net_2985), .C1(x3028) );
CLKBUF_X2 inst_9718 ( .A(net_9565), .Z(net_9566) );
SDFF_X2 inst_1543 ( .Q(net_7998), .D(net_7998), .SI(net_2712), .SE(net_2542), .CK(net_14414) );
CLKBUF_X2 inst_16954 ( .A(net_16801), .Z(net_16802) );
CLKBUF_X2 inst_16214 ( .A(net_15163), .Z(net_16062) );
CLKBUF_X2 inst_13892 ( .A(net_13739), .Z(net_13740) );
DFFR_X2 inst_7290 ( .QN(net_301), .D(net_300), .CK(net_16581), .RN(x6501) );
SDFF_X2 inst_1118 ( .D(net_7322), .SI(net_6564), .Q(net_6564), .SE(net_3070), .CK(net_11368) );
CLKBUF_X2 inst_15341 ( .A(net_15188), .Z(net_15189) );
DFFR_X2 inst_6978 ( .QN(net_5976), .D(net_5907), .CK(net_11553), .RN(x6501) );
INV_X4 inst_6109 ( .A(net_7494), .ZN(net_2968) );
CLKBUF_X2 inst_17768 ( .A(net_17615), .Z(net_17616) );
CLKBUF_X2 inst_10948 ( .A(net_10795), .Z(net_10796) );
SDFF_X2 inst_473 ( .SI(net_8479), .Q(net_8479), .SE(net_3983), .D(net_3939), .CK(net_12548) );
CLKBUF_X2 inst_15114 ( .A(net_14961), .Z(net_14962) );
CLKBUF_X2 inst_10140 ( .A(net_9987), .Z(net_9988) );
CLKBUF_X2 inst_16258 ( .A(net_16105), .Z(net_16106) );
CLKBUF_X2 inst_17303 ( .A(net_17150), .Z(net_17151) );
SDFFR_X2 inst_2211 ( .Q(net_7462), .D(net_7462), .SE(net_2863), .CK(net_10632), .SI(x13494), .RN(x6501) );
OAI21_X2 inst_3083 ( .B1(net_7635), .ZN(net_3155), .A(net_3154), .B2(net_3153) );
AND2_X2 inst_9170 ( .ZN(net_2505), .A2(net_2504), .A1(net_2391) );
CLKBUF_X2 inst_12609 ( .A(net_12456), .Z(net_12457) );
CLKBUF_X2 inst_15336 ( .A(net_15183), .Z(net_15184) );
CLKBUF_X2 inst_9917 ( .A(net_9764), .Z(net_9765) );
CLKBUF_X2 inst_12942 ( .A(net_12789), .Z(net_12790) );
CLKBUF_X2 inst_18821 ( .A(net_9586), .Z(net_18669) );
CLKBUF_X2 inst_15371 ( .A(net_15218), .Z(net_15219) );
CLKBUF_X2 inst_11034 ( .A(net_10881), .Z(net_10882) );
SDFF_X2 inst_1404 ( .SI(net_7277), .Q(net_7054), .D(net_7054), .SE(net_6280), .CK(net_17398) );
OAI21_X2 inst_2989 ( .ZN(net_5905), .B2(net_5902), .A(net_5821), .B1(net_691) );
INV_X4 inst_5880 ( .A(net_7604), .ZN(net_1760) );
NOR2_X2 inst_3479 ( .ZN(net_2405), .A1(net_2246), .A2(net_2245) );
NAND2_X2 inst_4704 ( .ZN(net_2715), .A1(net_1864), .A2(net_1586) );
NOR2_X2 inst_3575 ( .A1(net_7304), .ZN(net_1114), .A2(net_809) );
CLKBUF_X2 inst_9238 ( .A(net_9058), .Z(net_9086) );
NAND2_X2 inst_4493 ( .A1(net_7182), .A2(net_5655), .ZN(net_4479) );
AOI22_X2 inst_8484 ( .B1(net_6544), .A1(net_6511), .A2(net_6137), .B2(net_6104), .ZN(net_3456) );
CLKBUF_X2 inst_10180 ( .A(net_10027), .Z(net_10028) );
DFFR_X2 inst_7251 ( .QN(net_7305), .D(net_2045), .CK(net_15044), .RN(x6501) );
INV_X4 inst_5669 ( .A(net_8294), .ZN(net_956) );
CLKBUF_X2 inst_16556 ( .A(net_16403), .Z(net_16404) );
CLKBUF_X2 inst_10941 ( .A(net_10788), .Z(net_10789) );
SDFF_X2 inst_1395 ( .SI(net_7719), .Q(net_7719), .D(net_2576), .SE(net_2559), .CK(net_16064) );
SDFFR_X2 inst_2477 ( .Q(net_8986), .D(net_8986), .SI(net_2612), .SE(net_2562), .CK(net_14537), .RN(x6501) );
CLKBUF_X2 inst_14660 ( .A(net_14507), .Z(net_14508) );
INV_X4 inst_5460 ( .ZN(net_768), .A(net_767) );
CLKBUF_X2 inst_17316 ( .A(net_9141), .Z(net_17164) );
CLKBUF_X2 inst_11424 ( .A(net_11271), .Z(net_11272) );
AOI22_X2 inst_8322 ( .B1(net_8734), .A1(net_8512), .B2(net_4350), .A2(net_4349), .ZN(net_3724) );
NAND2_X2 inst_4838 ( .A1(net_7164), .ZN(net_1921), .A2(net_864) );
SDFF_X2 inst_1875 ( .D(net_7281), .SI(net_6978), .Q(net_6978), .SE(net_6283), .CK(net_18987) );
CLKBUF_X2 inst_10005 ( .A(net_9852), .Z(net_9853) );
OAI211_X2 inst_3190 ( .C2(net_7163), .C1(net_7162), .ZN(net_4725), .B(net_4417), .A(net_710) );
AOI22_X2 inst_8459 ( .B1(net_6605), .A1(net_6572), .A2(net_6257), .B2(net_6110), .ZN(net_3481) );
CLKBUF_X2 inst_10873 ( .A(net_9120), .Z(net_10721) );
NOR2_X2 inst_3397 ( .ZN(net_4515), .A1(net_4369), .A2(net_4368) );
CLKBUF_X2 inst_13286 ( .A(net_10514), .Z(net_13134) );
INV_X4 inst_5484 ( .A(net_959), .ZN(net_732) );
CLKBUF_X2 inst_11544 ( .A(net_11391), .Z(net_11392) );
NAND2_X2 inst_4421 ( .A1(net_6841), .A2(net_5016), .ZN(net_5006) );
AOI22_X2 inst_8448 ( .B1(net_6536), .A1(net_6503), .A2(net_6137), .B2(net_6104), .ZN(net_3492) );
NAND2_X2 inst_4233 ( .A1(net_6881), .A2(net_5247), .ZN(net_5227) );
DFFR_X2 inst_7128 ( .QN(net_7606), .D(net_3044), .CK(net_9782), .RN(x6501) );
INV_X4 inst_5905 ( .A(net_6389), .ZN(net_883) );
NAND3_X2 inst_3968 ( .ZN(net_2316), .A1(net_2315), .A3(net_2314), .A2(net_1932) );
CLKBUF_X2 inst_16535 ( .A(net_16382), .Z(net_16383) );
AOI22_X2 inst_8208 ( .B1(net_8867), .A1(net_8312), .B2(net_6252), .A2(net_4345), .ZN(net_3828) );
CLKBUF_X2 inst_19023 ( .A(net_13211), .Z(net_18871) );
CLKBUF_X2 inst_13010 ( .A(net_12857), .Z(net_12858) );
NAND2_X2 inst_4633 ( .ZN(net_2487), .A2(net_2443), .A1(net_2405) );
CLKBUF_X2 inst_16349 ( .A(net_16196), .Z(net_16197) );
AOI22_X2 inst_8113 ( .B1(net_7911), .A1(net_7809), .B2(net_6103), .A2(net_4398), .ZN(net_4035) );
CLKBUF_X2 inst_15845 ( .A(net_15692), .Z(net_15693) );
CLKBUF_X2 inst_14871 ( .A(net_13432), .Z(net_14719) );
HA_X1 inst_6660 ( .A(net_6174), .S(net_3987), .CO(net_3986), .B(net_1095) );
CLKBUF_X2 inst_10915 ( .A(net_10762), .Z(net_10763) );
AOI22_X2 inst_8027 ( .B1(net_8032), .A1(net_7998), .B2(net_6102), .A2(net_6097), .ZN(net_4110) );
INV_X2 inst_6411 ( .A(net_1151), .ZN(net_873) );
CLKBUF_X2 inst_9525 ( .A(net_9372), .Z(net_9373) );
AOI221_X2 inst_8769 ( .C1(net_8985), .B2(net_5538), .C2(net_5456), .ZN(net_5279), .A(net_4875), .B1(net_414) );
SDFF_X2 inst_618 ( .SI(net_8529), .Q(net_8529), .SE(net_3979), .D(net_3960), .CK(net_12270) );
SDFFR_X2 inst_2444 ( .SE(net_2685), .D(net_2667), .SI(net_471), .Q(net_471), .CK(net_16899), .RN(x6501) );
CLKBUF_X2 inst_11980 ( .A(net_11827), .Z(net_11828) );
OAI21_X2 inst_3057 ( .B2(net_8241), .B1(net_4850), .ZN(net_4750), .A(net_2597) );
SDFFR_X2 inst_2462 ( .SI(net_7377), .SE(net_2723), .D(net_2634), .QN(net_158), .CK(net_15035), .RN(x6501) );
HA_X1 inst_6706 ( .S(net_2177), .CO(net_1695), .A(net_1694), .B(net_1278) );
SDFF_X2 inst_474 ( .SI(net_8480), .Q(net_8480), .SE(net_3983), .D(net_3949), .CK(net_10577) );
CLKBUF_X2 inst_18865 ( .A(net_18712), .Z(net_18713) );
INV_X4 inst_5561 ( .A(net_1615), .ZN(net_608) );
SDFF_X2 inst_626 ( .SI(net_8520), .Q(net_8520), .SE(net_3979), .D(net_3943), .CK(net_13342) );
CLKBUF_X2 inst_15955 ( .A(net_15802), .Z(net_15803) );
CLKBUF_X2 inst_15560 ( .A(net_13287), .Z(net_15408) );
CLKBUF_X2 inst_14497 ( .A(net_12502), .Z(net_14345) );
CLKBUF_X2 inst_11539 ( .A(net_11386), .Z(net_11387) );
CLKBUF_X2 inst_9879 ( .A(net_9726), .Z(net_9727) );
DFFR_X1 inst_7476 ( .QN(net_7435), .D(net_3989), .CK(net_10115), .RN(x6501) );
CLKBUF_X2 inst_18143 ( .A(net_9539), .Z(net_17991) );
CLKBUF_X2 inst_16568 ( .A(net_13747), .Z(net_16416) );
CLKBUF_X2 inst_10247 ( .A(net_10094), .Z(net_10095) );
AOI21_X2 inst_8880 ( .B2(net_5871), .ZN(net_5864), .A(net_5863), .B1(x154) );
CLKBUF_X2 inst_11457 ( .A(net_10869), .Z(net_11305) );
CLKBUF_X2 inst_12641 ( .A(net_10811), .Z(net_12489) );
SDFF_X2 inst_798 ( .SI(net_8337), .Q(net_8337), .D(net_3977), .SE(net_3880), .CK(net_10712) );
CLKBUF_X2 inst_12648 ( .A(net_12495), .Z(net_12496) );
CLKBUF_X2 inst_16382 ( .A(net_16229), .Z(net_16230) );
CLKBUF_X2 inst_18215 ( .A(net_18062), .Z(net_18063) );
CLKBUF_X2 inst_16838 ( .A(net_16685), .Z(net_16686) );
NAND2_X2 inst_4340 ( .A1(net_7064), .A2(net_5162), .ZN(net_5117) );
SDFF_X2 inst_1434 ( .SI(net_7275), .Q(net_7092), .D(net_7092), .SE(net_6278), .CK(net_14641) );
CLKBUF_X2 inst_12727 ( .A(net_10966), .Z(net_12575) );
SDFF_X2 inst_1886 ( .D(net_7298), .SI(net_6995), .Q(net_6995), .SE(net_6283), .CK(net_18180) );
CLKBUF_X2 inst_18357 ( .A(net_18204), .Z(net_18205) );
CLKBUF_X2 inst_10211 ( .A(net_9643), .Z(net_10059) );
CLKBUF_X2 inst_16435 ( .A(net_16282), .Z(net_16283) );
CLKBUF_X2 inst_12889 ( .A(net_12736), .Z(net_12737) );
AOI221_X2 inst_8831 ( .C1(net_8147), .B1(net_7705), .C2(net_6101), .B2(net_6095), .ZN(net_6011), .A(net_4299) );
AOI221_X2 inst_8778 ( .C2(net_5535), .ZN(net_5261), .B2(net_5260), .A(net_4920), .B1(net_4890), .C1(net_448) );
NAND2_X2 inst_4349 ( .A1(net_7067), .A2(net_5162), .ZN(net_5108) );
SDFF_X2 inst_1457 ( .SI(net_7275), .Q(net_7132), .D(net_7132), .SE(net_6279), .CK(net_17385) );
AOI222_X1 inst_8627 ( .A2(net_8219), .C2(net_6117), .A1(net_4800), .B2(net_4799), .ZN(net_4797), .B1(net_3138), .C1(net_2101) );
CLKBUF_X2 inst_10552 ( .A(net_9706), .Z(net_10400) );
CLKBUF_X2 inst_16635 ( .A(net_16482), .Z(net_16483) );
CLKBUF_X2 inst_13244 ( .A(net_13091), .Z(net_13092) );
AOI22_X2 inst_8209 ( .B1(net_8831), .A1(net_8350), .A2(net_6265), .B2(net_6253), .ZN(net_3827) );
CLKBUF_X2 inst_11254 ( .A(net_11101), .Z(net_11102) );
NAND4_X2 inst_3662 ( .A4(net_6014), .A1(net_6013), .ZN(net_4603), .A2(net_4120), .A3(net_4119) );
CLKBUF_X2 inst_18117 ( .A(net_17964), .Z(net_17965) );
SDFFR_X1 inst_2670 ( .D(net_6785), .SE(net_4506), .CK(net_11407), .RN(x6501), .SI(x1281), .Q(x1281) );
CLKBUF_X2 inst_15726 ( .A(net_15573), .Z(net_15574) );
CLKBUF_X2 inst_10983 ( .A(net_10723), .Z(net_10831) );
AOI22_X2 inst_8380 ( .B1(net_8671), .A1(net_8634), .B2(net_6109), .A2(net_3857), .ZN(net_3668) );
OAI221_X2 inst_2974 ( .A(net_2433), .ZN(net_2431), .B1(net_2277), .B2(net_831), .C1(net_731), .C2(net_635) );
CLKBUF_X2 inst_16965 ( .A(net_16812), .Z(net_16813) );
SDFF_X2 inst_1895 ( .D(net_7285), .SI(net_7022), .Q(net_7022), .SE(net_6277), .CK(net_16183) );
AOI22_X2 inst_8476 ( .B1(net_6542), .A1(net_6509), .A2(net_6137), .B2(net_6104), .ZN(net_3464) );
SDFFR_X1 inst_2730 ( .SI(net_9043), .Q(net_9043), .D(net_7472), .SE(net_3208), .CK(net_12213), .RN(x6501) );
CLKBUF_X2 inst_19159 ( .A(net_19006), .Z(net_19007) );
SDFF_X2 inst_737 ( .SI(net_8352), .Q(net_8352), .D(net_3958), .SE(net_3880), .CK(net_9996) );
CLKBUF_X2 inst_11725 ( .A(net_11572), .Z(net_11573) );
CLKBUF_X2 inst_11178 ( .A(net_11025), .Z(net_11026) );
CLKBUF_X2 inst_16373 ( .A(net_11144), .Z(net_16221) );
AOI21_X2 inst_8990 ( .B1(net_5953), .ZN(net_3939), .A(net_1458), .B2(net_1054) );
SDFF_X2 inst_545 ( .Q(net_8689), .D(net_8689), .SI(net_3963), .SE(net_3935), .CK(net_10070) );
CLKBUF_X2 inst_16905 ( .A(net_16752), .Z(net_16753) );
CLKBUF_X2 inst_15819 ( .A(net_15666), .Z(net_15667) );
AOI22_X2 inst_8373 ( .B1(net_8670), .A1(net_8633), .B2(net_6109), .A2(net_3857), .ZN(net_3675) );
CLKBUF_X2 inst_10189 ( .A(net_9466), .Z(net_10037) );
AOI22_X2 inst_8132 ( .B1(net_8185), .A1(net_7675), .B2(net_6099), .A2(net_4399), .ZN(net_4017) );
CLKBUF_X2 inst_17733 ( .A(net_15747), .Z(net_17581) );
DFF_X1 inst_6854 ( .Q(net_6442), .D(net_3627), .CK(net_17891) );
CLKBUF_X2 inst_14475 ( .A(net_14322), .Z(net_14323) );
CLKBUF_X2 inst_12188 ( .A(net_12035), .Z(net_12036) );
HA_X1 inst_6682 ( .A(net_3236), .S(net_3041), .CO(net_3040), .B(net_2872) );
CLKBUF_X2 inst_13595 ( .A(net_13442), .Z(net_13443) );
AOI22_X2 inst_7832 ( .A2(net_5535), .B2(net_5260), .ZN(net_4689), .B1(net_3309), .A1(net_456) );
AOI222_X1 inst_8624 ( .A2(net_8252), .B1(net_7594), .C2(net_6116), .ZN(net_4802), .A1(net_4800), .B2(net_4799), .C1(net_2571) );
INV_X4 inst_5878 ( .A(net_6397), .ZN(net_2754) );
CLKBUF_X2 inst_14383 ( .A(net_14230), .Z(net_14231) );
AOI21_X2 inst_8910 ( .ZN(net_5790), .A(net_5746), .B2(net_5656), .B1(net_4911) );
CLKBUF_X2 inst_13356 ( .A(net_13091), .Z(net_13204) );
INV_X2 inst_6573 ( .ZN(net_799), .A(net_217) );
CLKBUF_X2 inst_13067 ( .A(net_12914), .Z(net_12915) );
CLKBUF_X2 inst_12347 ( .A(net_12194), .Z(net_12195) );
CLKBUF_X2 inst_10559 ( .A(net_9516), .Z(net_10407) );
CLKBUF_X2 inst_13879 ( .A(net_13369), .Z(net_13727) );
NAND2_X2 inst_4415 ( .A1(net_6854), .A2(net_5016), .ZN(net_5012) );
NAND2_X2 inst_4209 ( .ZN(net_5271), .A2(net_5270), .A1(net_2207) );
CLKBUF_X2 inst_10266 ( .A(net_9271), .Z(net_10114) );
INV_X16 inst_6635 ( .ZN(net_3969), .A(net_3360) );
CLKBUF_X2 inst_15932 ( .A(net_15779), .Z(net_15780) );
CLKBUF_X2 inst_10275 ( .A(net_9755), .Z(net_10123) );
CLKBUF_X2 inst_18746 ( .A(net_18593), .Z(net_18594) );
AOI22_X2 inst_8561 ( .A1(net_2634), .ZN(net_2335), .A2(net_2334), .B2(net_2333), .B1(net_1757) );
AOI21_X2 inst_8972 ( .B2(net_5950), .A(net_2483), .ZN(net_2476), .B1(net_918) );
CLKBUF_X2 inst_16781 ( .A(net_16628), .Z(net_16629) );
CLKBUF_X2 inst_12072 ( .A(net_11919), .Z(net_11920) );
INV_X4 inst_5828 ( .A(net_6305), .ZN(net_2686) );
NAND2_X2 inst_4260 ( .A1(net_7032), .A2(net_5249), .ZN(net_5200) );
CLKBUF_X2 inst_10218 ( .A(net_9534), .Z(net_10066) );
AOI22_X2 inst_8072 ( .B1(net_7937), .A1(net_7835), .B2(net_6103), .A2(net_4398), .ZN(net_4072) );
NOR2_X2 inst_3484 ( .A1(net_3023), .ZN(net_2226), .A2(net_2032) );
CLKBUF_X2 inst_13868 ( .A(net_13715), .Z(net_13716) );
SDFF_X2 inst_942 ( .SI(net_7323), .Q(net_6697), .D(net_6697), .SE(net_3125), .CK(net_9147) );
AOI22_X2 inst_7755 ( .B1(net_6983), .A1(net_6943), .A2(net_5443), .B2(net_5442), .ZN(net_5386) );
CLKBUF_X2 inst_12077 ( .A(net_11924), .Z(net_11925) );
AOI22_X2 inst_8269 ( .B1(net_8875), .A1(net_8320), .B2(net_6252), .A2(net_4345), .ZN(net_3769) );
CLKBUF_X2 inst_13174 ( .A(net_13021), .Z(net_13022) );
INV_X2 inst_6603 ( .A(net_6161), .ZN(net_6160) );
DFFR_X2 inst_7338 ( .Q(net_7339), .CK(net_11719), .D(x12922), .RN(x6501) );
DFFR_X2 inst_7353 ( .Q(net_7312), .CK(net_11375), .D(x13174), .RN(x6501) );
NAND2_X2 inst_4501 ( .ZN(net_4386), .A1(net_4385), .A2(net_4319) );
DFFR_X2 inst_7144 ( .QN(net_7518), .D(net_2884), .CK(net_14829), .RN(x6501) );
NAND2_X2 inst_4252 ( .A1(net_7029), .A2(net_5249), .ZN(net_5208) );
CLKBUF_X2 inst_11758 ( .A(net_10815), .Z(net_11606) );
INV_X2 inst_6356 ( .ZN(net_2197), .A(net_2196) );
AOI22_X2 inst_8258 ( .B1(net_8763), .A1(net_8393), .A2(net_3867), .B2(net_3866), .ZN(net_3780) );
CLKBUF_X2 inst_18728 ( .A(net_11149), .Z(net_18576) );
INV_X4 inst_5451 ( .ZN(net_1427), .A(net_805) );
CLKBUF_X2 inst_16929 ( .A(net_16776), .Z(net_16777) );
CLKBUF_X2 inst_16124 ( .A(net_15971), .Z(net_15972) );
INV_X2 inst_6393 ( .ZN(net_1179), .A(net_1178) );
SDFF_X2 inst_418 ( .SI(net_8333), .Q(net_8333), .SE(net_3978), .D(net_3948), .CK(net_13488) );
CLKBUF_X2 inst_17368 ( .A(net_17215), .Z(net_17216) );
NAND3_X2 inst_3961 ( .ZN(net_4774), .A1(net_2843), .A2(net_2764), .A3(net_2642) );
CLKBUF_X2 inst_19155 ( .A(net_19002), .Z(net_19003) );
CLKBUF_X2 inst_9526 ( .A(net_9373), .Z(net_9374) );
CLKBUF_X2 inst_11851 ( .A(net_11698), .Z(net_11699) );
INV_X4 inst_5871 ( .A(net_8935), .ZN(net_2602) );
CLKBUF_X2 inst_10016 ( .A(net_9505), .Z(net_9864) );
CLKBUF_X2 inst_16241 ( .A(net_16088), .Z(net_16089) );
CLKBUF_X2 inst_13957 ( .A(net_13804), .Z(net_13805) );
SDFF_X2 inst_1177 ( .SI(net_7315), .Q(net_6590), .D(net_6590), .SE(net_3069), .CK(net_9895) );
SDFFR_X2 inst_2548 ( .QN(net_6359), .SE(net_2147), .D(net_2136), .SI(net_1952), .CK(net_17405), .RN(x6501) );
CLKBUF_X2 inst_11494 ( .A(net_11341), .Z(net_11342) );
INV_X4 inst_5127 ( .ZN(net_4486), .A(net_4382) );
AOI22_X2 inst_8022 ( .A1(net_7964), .B1(net_7794), .A2(net_6092), .B2(net_6091), .ZN(net_4114) );
CLKBUF_X2 inst_12587 ( .A(net_12434), .Z(net_12435) );
AND3_X2 inst_9051 ( .A3(net_2123), .A1(net_1284), .A2(net_1280), .ZN(net_1056) );
SDFF_X2 inst_1666 ( .SI(net_7762), .Q(net_7762), .D(net_2717), .SE(net_2560), .CK(net_13762) );
CLKBUF_X2 inst_17916 ( .A(net_17763), .Z(net_17764) );
SDFF_X2 inst_735 ( .SI(net_8348), .Q(net_8348), .D(net_3959), .SE(net_3880), .CK(net_13186) );
SDFF_X2 inst_1529 ( .Q(net_7906), .D(net_7906), .SI(net_2656), .SE(net_2543), .CK(net_16723) );
CLKBUF_X2 inst_18992 ( .A(net_18839), .Z(net_18840) );
CLKBUF_X2 inst_16798 ( .A(net_11178), .Z(net_16646) );
CLKBUF_X2 inst_12445 ( .A(net_12292), .Z(net_12293) );
CLKBUF_X2 inst_10426 ( .A(net_10273), .Z(net_10274) );
AOI22_X2 inst_7890 ( .A2(net_4809), .ZN(net_4541), .B1(net_4540), .B2(net_4388), .A1(net_347) );
SDFF_X2 inst_1653 ( .SI(net_7737), .Q(net_7737), .D(net_2703), .SE(net_2559), .CK(net_14004) );
CLKBUF_X2 inst_17230 ( .A(net_17077), .Z(net_17078) );
CLKBUF_X2 inst_18777 ( .A(net_18624), .Z(net_18625) );
CLKBUF_X2 inst_13376 ( .A(net_13223), .Z(net_13224) );
DFFR_X2 inst_7220 ( .D(net_2369), .QN(net_214), .CK(net_17878), .RN(x6501) );
CLKBUF_X2 inst_18052 ( .A(net_17899), .Z(net_17900) );
CLKBUF_X2 inst_11627 ( .A(net_11474), .Z(net_11475) );
OAI21_X2 inst_2984 ( .ZN(net_5926), .A(net_5851), .B2(net_3060), .B1(net_2460) );
NOR3_X2 inst_3258 ( .ZN(net_4501), .A3(net_4390), .A1(net_4325), .A2(net_1347) );
CLKBUF_X2 inst_13002 ( .A(net_12849), .Z(net_12850) );
CLKBUF_X2 inst_12150 ( .A(net_11690), .Z(net_11998) );
SDFF_X2 inst_1805 ( .D(net_7270), .SI(net_6927), .Q(net_6927), .SE(net_6281), .CK(net_14355) );
NOR2_X2 inst_3563 ( .A1(net_7364), .ZN(net_1293), .A2(net_1292) );
CLKBUF_X2 inst_18339 ( .A(net_10868), .Z(net_18187) );
CLKBUF_X2 inst_16628 ( .A(net_16475), .Z(net_16476) );
CLKBUF_X2 inst_9675 ( .A(net_9522), .Z(net_9523) );
CLKBUF_X2 inst_16088 ( .A(net_15935), .Z(net_15936) );
AOI22_X2 inst_8231 ( .B1(net_8760), .A1(net_8390), .A2(net_3867), .B2(net_3866), .ZN(net_3806) );
AOI21_X2 inst_8936 ( .B2(net_5871), .ZN(net_5667), .A(net_5666), .B1(net_2687) );
SDFFR_X1 inst_2752 ( .QN(net_7561), .D(net_3961), .SI(net_3145), .SE(net_3144), .CK(net_11036), .RN(x6501) );
CLKBUF_X2 inst_10095 ( .A(net_9942), .Z(net_9943) );
CLKBUF_X2 inst_16140 ( .A(net_15987), .Z(net_15988) );
SDFF_X2 inst_1281 ( .Q(net_8081), .D(net_8081), .SE(net_2707), .SI(net_2655), .CK(net_15549) );
CLKBUF_X2 inst_19032 ( .A(net_18879), .Z(net_18880) );
SDFF_X2 inst_1509 ( .SI(net_7842), .Q(net_7842), .D(net_2705), .SE(net_2558), .CK(net_18551) );
OAI21_X2 inst_3088 ( .ZN(net_2948), .B2(net_2947), .B1(net_2945), .A(net_2906) );
CLKBUF_X2 inst_10386 ( .A(net_10233), .Z(net_10234) );
AOI21_X2 inst_9000 ( .A(net_1333), .ZN(net_1272), .B1(net_1271), .B2(net_909) );
CLKBUF_X2 inst_15858 ( .A(net_15705), .Z(net_15706) );
NAND4_X2 inst_3782 ( .ZN(net_4239), .A1(net_3691), .A2(net_3690), .A3(net_3689), .A4(net_3688) );
CLKBUF_X2 inst_15754 ( .A(net_15601), .Z(net_15602) );
DFFR_X1 inst_7486 ( .QN(net_7422), .D(net_4228), .CK(net_12311), .RN(x6501) );
CLKBUF_X2 inst_15101 ( .A(net_10528), .Z(net_14949) );
CLKBUF_X2 inst_15466 ( .A(net_15313), .Z(net_15314) );
INV_X16 inst_6630 ( .ZN(net_4350), .A(net_3377) );
CLKBUF_X2 inst_15378 ( .A(net_15225), .Z(net_15226) );
AOI22_X2 inst_8054 ( .B1(net_8104), .A1(net_7764), .B2(net_6108), .A2(net_6096), .ZN(net_4087) );
INV_X4 inst_5809 ( .A(net_8279), .ZN(net_680) );
SDFF_X2 inst_1140 ( .D(net_7319), .SI(net_6561), .Q(net_6561), .SE(net_3070), .CK(net_9840) );
CLKBUF_X2 inst_15637 ( .A(net_15484), .Z(net_15485) );
CLKBUF_X2 inst_9251 ( .A(net_9098), .Z(net_9099) );
INV_X4 inst_6140 ( .A(net_6118), .ZN(net_6117) );
SDFF_X2 inst_1800 ( .D(net_7274), .SI(net_6971), .Q(net_6971), .SE(net_6283), .CK(net_17376) );
NAND2_X2 inst_4773 ( .ZN(net_2401), .A2(net_2307), .A1(net_1639) );
AOI22_X2 inst_8463 ( .B1(net_6521), .A1(net_6488), .A2(net_6137), .B2(net_6104), .ZN(net_3477) );
CLKBUF_X2 inst_11087 ( .A(net_10934), .Z(net_10935) );
SDFF_X2 inst_448 ( .Q(net_8745), .D(net_8745), .SE(net_3982), .SI(net_3938), .CK(net_13060) );
INV_X4 inst_5966 ( .A(net_6460), .ZN(net_516) );
INV_X4 inst_5680 ( .A(net_7663), .ZN(net_1553) );
CLKBUF_X2 inst_10253 ( .A(net_10100), .Z(net_10101) );
INV_X4 inst_6056 ( .A(net_5968), .ZN(x3207) );
MUX2_X2 inst_4921 ( .B(net_6817), .S(net_6272), .Z(net_4620), .A(net_4619) );
CLKBUF_X2 inst_14367 ( .A(net_14214), .Z(net_14215) );
CLKBUF_X2 inst_9374 ( .A(net_9177), .Z(net_9222) );
CLKBUF_X2 inst_10862 ( .A(net_10709), .Z(net_10710) );
CLKBUF_X2 inst_10053 ( .A(net_9440), .Z(net_9901) );
CLKBUF_X2 inst_16072 ( .A(net_15919), .Z(net_15920) );
CLKBUF_X2 inst_18624 ( .A(net_18471), .Z(net_18472) );
CLKBUF_X2 inst_13017 ( .A(net_11729), .Z(net_12865) );
AOI22_X2 inst_8212 ( .B1(net_8794), .A1(net_8535), .A2(net_3861), .B2(net_3860), .ZN(net_3824) );
SDFF_X2 inst_1343 ( .Q(net_8181), .D(net_8181), .SI(net_2585), .SE(net_2561), .CK(net_18563) );
AND2_X4 inst_9068 ( .A1(net_6169), .ZN(net_5043), .A2(net_3217) );
AOI22_X2 inst_8050 ( .B1(net_8138), .A1(net_7900), .A2(net_6098), .ZN(net_6042), .B2(net_4190) );
CLKBUF_X2 inst_16133 ( .A(net_15980), .Z(net_15981) );
DFFR_X1 inst_7536 ( .Q(net_7170), .D(net_590), .CK(net_11847), .RN(x6501) );
NAND2_X4 inst_4054 ( .A2(net_7210), .ZN(net_1802), .A1(net_692) );
AOI22_X2 inst_7813 ( .A2(net_8246), .B2(net_6144), .A1(net_4764), .ZN(net_4745), .B1(net_4540) );
HA_X1 inst_6713 ( .B(net_2997), .A(net_2989), .S(net_1231), .CO(net_1230) );
SDFF_X2 inst_1246 ( .SI(net_7690), .Q(net_7690), .D(net_2718), .SE(net_2714), .CK(net_18819) );
OAI211_X2 inst_3185 ( .ZN(net_5523), .C2(net_5036), .B(net_4730), .A(net_1519), .C1(net_1161) );
CLKBUF_X2 inst_17419 ( .A(net_16527), .Z(net_17267) );
NAND2_X2 inst_4679 ( .A2(net_2299), .ZN(net_2253), .A1(net_2089) );
CLKBUF_X2 inst_11699 ( .A(net_9346), .Z(net_11547) );
CLKBUF_X2 inst_11269 ( .A(net_11116), .Z(net_11117) );
CLKBUF_X2 inst_13163 ( .A(net_13010), .Z(net_13011) );
CLKBUF_X2 inst_15881 ( .A(net_15728), .Z(net_15729) );
INV_X4 inst_5647 ( .A(net_6834), .ZN(net_2104) );
CLKBUF_X2 inst_10623 ( .A(net_10470), .Z(net_10471) );
INV_X4 inst_5580 ( .A(net_9005), .ZN(net_2529) );
CLKBUF_X2 inst_12180 ( .A(net_12027), .Z(net_12028) );
CLKBUF_X2 inst_16351 ( .A(net_16198), .Z(net_16199) );
AOI22_X2 inst_8568 ( .ZN(net_2165), .A1(net_2164), .B2(net_2163), .A2(net_2082), .B1(net_2081) );
SDFF_X2 inst_2029 ( .SI(net_7935), .Q(net_7935), .D(net_2639), .SE(net_2461), .CK(net_16450) );
CLKBUF_X2 inst_17298 ( .A(net_17145), .Z(net_17146) );
CLKBUF_X2 inst_10632 ( .A(net_10195), .Z(net_10480) );
CLKBUF_X2 inst_12812 ( .A(net_12659), .Z(net_12660) );
AOI221_X2 inst_8779 ( .C2(net_5535), .B2(net_5260), .ZN(net_5259), .A(net_4919), .B1(net_4884), .C1(net_451) );
MUX2_X2 inst_4936 ( .B(net_8964), .A(net_3003), .S(net_2967), .Z(net_2890) );
CLKBUF_X2 inst_15037 ( .A(net_14884), .Z(net_14885) );
CLKBUF_X2 inst_16528 ( .A(net_16375), .Z(net_16376) );
CLKBUF_X2 inst_18784 ( .A(net_18631), .Z(net_18632) );
SDFF_X2 inst_1965 ( .D(net_7271), .SI(net_6848), .Q(net_6848), .SE(net_6282), .CK(net_14074) );
CLKBUF_X2 inst_16033 ( .A(net_15880), .Z(net_15881) );
NAND3_X2 inst_3915 ( .ZN(net_5623), .A1(net_5552), .A3(net_5486), .A2(net_5333) );
INV_X4 inst_5419 ( .A(net_1267), .ZN(net_859) );
AOI22_X2 inst_8144 ( .B1(net_7915), .A1(net_7813), .B2(net_6103), .A2(net_4398), .ZN(net_4007) );
INV_X4 inst_5743 ( .A(net_7420), .ZN(net_2150) );
CLKBUF_X2 inst_19127 ( .A(net_18974), .Z(net_18975) );
INV_X4 inst_5422 ( .ZN(net_2530), .A(net_856) );
CLKBUF_X2 inst_18913 ( .A(net_18760), .Z(net_18761) );
CLKBUF_X2 inst_15785 ( .A(net_15064), .Z(net_15633) );
NOR3_X2 inst_3285 ( .ZN(net_2740), .A1(net_2400), .A2(net_2318), .A3(net_2317) );
DFFS_X1 inst_6948 ( .D(net_6145), .CK(net_13626), .SN(x6501), .Q(x712) );
INV_X2 inst_6492 ( .A(net_7356), .ZN(net_833) );
CLKBUF_X2 inst_14091 ( .A(net_13938), .Z(net_13939) );
CLKBUF_X2 inst_14934 ( .A(net_14395), .Z(net_14782) );
CLKBUF_X2 inst_11931 ( .A(net_11778), .Z(net_11779) );
CLKBUF_X2 inst_11790 ( .A(net_11469), .Z(net_11638) );
CLKBUF_X2 inst_11568 ( .A(net_11415), .Z(net_11416) );
NAND2_X2 inst_4460 ( .ZN(net_4932), .A2(net_4711), .A1(net_4493) );
CLKBUF_X2 inst_18046 ( .A(net_14003), .Z(net_17894) );
AOI22_X2 inst_8336 ( .B1(net_8736), .A1(net_8514), .B2(net_4350), .A2(net_4349), .ZN(net_3711) );
CLKBUF_X2 inst_12559 ( .A(net_12406), .Z(net_12407) );
CLKBUF_X2 inst_11681 ( .A(net_11528), .Z(net_11529) );
DFFR_X2 inst_7002 ( .D(net_5880), .CK(net_11435), .RN(x6501), .Q(x2542) );
OR3_X4 inst_2804 ( .ZN(net_1925), .A2(net_1057), .A1(x12843), .A3(x12780) );
INV_X4 inst_5131 ( .ZN(net_4555), .A(net_4368) );
SDFF_X2 inst_772 ( .Q(net_8783), .D(net_8783), .SI(net_3965), .SE(net_3879), .CK(net_12429) );
DFF_X1 inst_6738 ( .Q(net_6783), .D(net_5631), .CK(net_11426) );
NAND4_X2 inst_3682 ( .A4(net_6054), .A1(net_6053), .ZN(net_4583), .A2(net_3998), .A3(net_3997) );
MUX2_X2 inst_4940 ( .A(net_4671), .Z(net_2761), .B(net_2760), .S(net_2417) );
NAND2_X2 inst_4583 ( .A2(net_3033), .ZN(net_2950), .A1(net_2949) );
CLKBUF_X2 inst_13282 ( .A(net_12022), .Z(net_13130) );
CLKBUF_X2 inst_15141 ( .A(net_14335), .Z(net_14989) );
CLKBUF_X2 inst_10525 ( .A(net_10372), .Z(net_10373) );
CLKBUF_X2 inst_14396 ( .A(net_12641), .Z(net_14244) );
NAND2_X2 inst_4870 ( .ZN(net_2019), .A1(net_1316), .A2(net_827) );
INV_X4 inst_5454 ( .A(net_7210), .ZN(net_1481) );
CLKBUF_X2 inst_17047 ( .A(net_16367), .Z(net_16895) );
INV_X2 inst_6224 ( .ZN(net_5486), .A(net_5332) );
DFF_X1 inst_6761 ( .Q(net_7541), .D(net_4611), .CK(net_11971) );
SDFF_X2 inst_606 ( .SI(net_8373), .Q(net_8373), .D(net_3980), .SE(net_3969), .CK(net_13121) );
OAI22_X2 inst_2942 ( .A1(net_2097), .ZN(net_1878), .B1(net_1877), .A2(net_1613), .B2(net_1327) );
CLKBUF_X2 inst_9929 ( .A(net_9776), .Z(net_9777) );
CLKBUF_X2 inst_16496 ( .A(net_12889), .Z(net_16344) );
CLKBUF_X2 inst_13875 ( .A(net_10669), .Z(net_13723) );
CLKBUF_X2 inst_10287 ( .A(net_10134), .Z(net_10135) );
AOI22_X2 inst_8167 ( .B1(net_8825), .A1(net_8344), .A2(net_6265), .B2(net_6253), .ZN(net_3869) );
XNOR2_X2 inst_139 ( .A(net_6188), .ZN(net_2460), .B(x3327) );
CLKBUF_X2 inst_13767 ( .A(net_13614), .Z(net_13615) );
CLKBUF_X2 inst_15813 ( .A(net_15660), .Z(net_15661) );
CLKBUF_X2 inst_10856 ( .A(net_10703), .Z(net_10704) );
AOI21_X2 inst_8903 ( .B2(net_5871), .ZN(net_5763), .A(net_5762), .B1(net_2681) );
CLKBUF_X2 inst_12548 ( .A(net_9391), .Z(net_12396) );
SDFF_X2 inst_1316 ( .SI(net_7673), .Q(net_7673), .SE(net_2714), .D(net_2655), .CK(net_18571) );
AOI22_X2 inst_8400 ( .B1(net_8748), .A1(net_8378), .A2(net_3867), .B2(net_3866), .ZN(net_3652) );
NOR2_X2 inst_3551 ( .A1(net_1910), .ZN(net_1664), .A2(net_1591) );
INV_X4 inst_5528 ( .ZN(net_1043), .A(net_662) );
CLKBUF_X2 inst_18504 ( .A(net_12578), .Z(net_18352) );
INV_X2 inst_6521 ( .ZN(net_788), .A(net_223) );
XNOR2_X2 inst_191 ( .ZN(net_1572), .A(net_942), .B(net_937) );
CLKBUF_X2 inst_16552 ( .A(net_16399), .Z(net_16400) );
AOI21_X2 inst_8908 ( .ZN(net_5785), .A(net_5746), .B2(net_5652), .B1(net_4487) );
CLKBUF_X2 inst_9328 ( .A(net_9175), .Z(net_9176) );
CLKBUF_X2 inst_13485 ( .A(net_13332), .Z(net_13333) );
NAND2_X2 inst_4538 ( .A1(net_3371), .ZN(net_3370), .A2(net_3369) );
INV_X4 inst_5212 ( .ZN(net_2354), .A(net_2294) );
CLKBUF_X2 inst_13988 ( .A(net_13835), .Z(net_13836) );
CLKBUF_X2 inst_18279 ( .A(net_15743), .Z(net_18127) );
DFFS_X2 inst_6892 ( .QN(net_7356), .D(net_2855), .CK(net_11801), .SN(x6501) );
NAND3_X4 inst_3879 ( .ZN(net_6157), .A1(net_1630), .A3(net_1249), .A2(net_1248) );
INV_X4 inst_5269 ( .A(net_4956), .ZN(net_4685) );
CLKBUF_X2 inst_19143 ( .A(net_18990), .Z(net_18991) );
INV_X2 inst_6544 ( .A(net_6372), .ZN(net_2135) );
CLKBUF_X2 inst_12201 ( .A(net_12048), .Z(net_12049) );
SDFFR_X2 inst_2184 ( .SI(net_8894), .Q(net_8894), .SE(net_3022), .D(net_1424), .CK(net_18916), .RN(x6501) );
CLKBUF_X2 inst_13296 ( .A(net_13143), .Z(net_13144) );
SDFFR_X1 inst_2665 ( .D(net_6762), .SE(net_4506), .CK(net_11535), .RN(x6501), .SI(x2006), .Q(x2006) );
SDFF_X2 inst_1132 ( .D(net_7340), .SI(net_6582), .Q(net_6582), .SE(net_3070), .CK(net_9609) );
CLKBUF_X2 inst_14415 ( .A(net_14140), .Z(net_14263) );
CLKBUF_X2 inst_17619 ( .A(net_17466), .Z(net_17467) );
SDFF_X2 inst_968 ( .SI(net_7329), .Q(net_6736), .D(net_6736), .SE(net_3124), .CK(net_11650) );
NAND2_X2 inst_4700 ( .ZN(net_1873), .A1(net_1872), .A2(net_1871) );
CLKBUF_X2 inst_13531 ( .A(net_11899), .Z(net_13379) );
NAND2_X2 inst_4441 ( .A1(net_6878), .A2(net_5016), .ZN(net_4986) );
CLKBUF_X2 inst_15024 ( .A(net_13741), .Z(net_14872) );
OAI21_X2 inst_3153 ( .B2(net_1984), .ZN(net_1981), .A(net_1979), .B1(net_653) );
INV_X4 inst_6076 ( .A(net_5970), .ZN(x3288) );
CLKBUF_X2 inst_14357 ( .A(net_14204), .Z(net_14205) );
CLKBUF_X2 inst_11990 ( .A(net_11837), .Z(net_11838) );
NAND3_X2 inst_4004 ( .A3(net_1324), .A2(net_1322), .ZN(net_1301), .A1(net_619) );
CLKBUF_X2 inst_12708 ( .A(net_11075), .Z(net_12556) );
CLKBUF_X2 inst_15352 ( .A(net_15199), .Z(net_15200) );
CLKBUF_X2 inst_18513 ( .A(net_18360), .Z(net_18361) );
CLKBUF_X2 inst_17312 ( .A(net_17159), .Z(net_17160) );
CLKBUF_X2 inst_11838 ( .A(net_9347), .Z(net_11686) );
AOI21_X2 inst_8887 ( .B2(net_5871), .ZN(net_5811), .A(net_5805), .B1(x406) );
NAND4_X2 inst_3798 ( .ZN(net_3628), .A2(net_3500), .A1(net_3499), .A3(net_3498), .A4(net_3497) );
CLKBUF_X2 inst_18137 ( .A(net_17984), .Z(net_17985) );
INV_X4 inst_5232 ( .ZN(net_2418), .A(net_2165) );
NAND2_X2 inst_4109 ( .ZN(net_5421), .A1(net_5237), .A2(net_5011) );
NAND2_X2 inst_4192 ( .ZN(net_5308), .A2(net_5182), .A1(net_5063) );
CLKBUF_X2 inst_10048 ( .A(net_9291), .Z(net_9896) );
OAI21_X2 inst_3004 ( .ZN(net_5927), .B2(net_5739), .A(net_5718), .B1(net_4949) );
CLKBUF_X2 inst_12396 ( .A(net_12243), .Z(net_12244) );
NAND2_X2 inst_4672 ( .ZN(net_2370), .A2(net_2116), .A1(net_2115) );
CLKBUF_X2 inst_14438 ( .A(net_14285), .Z(net_14286) );
CLKBUF_X2 inst_12363 ( .A(net_12210), .Z(net_12211) );
CLKBUF_X2 inst_17355 ( .A(net_17202), .Z(net_17203) );
CLKBUF_X2 inst_17024 ( .A(net_16871), .Z(net_16872) );
SDFFR_X2 inst_2456 ( .SE(net_2354), .D(net_2293), .SI(net_269), .Q(net_269), .CK(net_16103), .RN(x6501) );
OR2_X2 inst_2887 ( .ZN(net_2010), .A2(net_1740), .A1(net_1669) );
CLKBUF_X2 inst_12162 ( .A(net_12009), .Z(net_12010) );
CLKBUF_X2 inst_11120 ( .A(net_10967), .Z(net_10968) );
CLKBUF_X2 inst_18655 ( .A(net_18502), .Z(net_18503) );
CLKBUF_X2 inst_16972 ( .A(net_16819), .Z(net_16820) );
AOI221_X2 inst_8805 ( .B1(net_7185), .C2(net_5657), .B2(net_5655), .A(net_4834), .ZN(net_4824), .C1(net_2634) );
SDFF_X2 inst_1473 ( .SI(net_7267), .Q(net_7124), .D(net_7124), .SE(net_6279), .CK(net_16845) );
INV_X4 inst_5334 ( .ZN(net_1478), .A(net_1467) );
CLKBUF_X2 inst_12793 ( .A(net_9156), .Z(net_12641) );
CLKBUF_X2 inst_9306 ( .A(net_9059), .Z(net_9154) );
CLKBUF_X2 inst_16248 ( .A(net_16095), .Z(net_16096) );
CLKBUF_X2 inst_18099 ( .A(net_17946), .Z(net_17947) );
SDFF_X2 inst_632 ( .SI(net_8546), .Q(net_8546), .SE(net_3979), .D(net_3941), .CK(net_12886) );
CLKBUF_X2 inst_18435 ( .A(net_18282), .Z(net_18283) );
XOR2_X2 inst_0 ( .B(net_7441), .Z(net_4314), .A(net_3986) );
CLKBUF_X2 inst_13934 ( .A(net_13781), .Z(net_13782) );
CLKBUF_X2 inst_17242 ( .A(net_17089), .Z(net_17090) );
CLKBUF_X2 inst_11405 ( .A(net_11252), .Z(net_11253) );
CLKBUF_X2 inst_14582 ( .A(net_14429), .Z(net_14430) );
CLKBUF_X2 inst_11199 ( .A(net_11046), .Z(net_11047) );
CLKBUF_X2 inst_12266 ( .A(net_12113), .Z(net_12114) );
AOI21_X2 inst_8994 ( .B2(net_1745), .ZN(net_1437), .A(net_1018), .B1(net_188) );
CLKBUF_X2 inst_13520 ( .A(net_9850), .Z(net_13368) );
SDFF_X2 inst_1983 ( .D(net_7275), .SI(net_6892), .Q(net_6892), .SE(net_6284), .CK(net_14598) );
CLKBUF_X2 inst_13748 ( .A(net_13595), .Z(net_13596) );
DFFR_X2 inst_7323 ( .QN(net_389), .D(net_297), .CK(net_18942), .RN(x6501) );
CLKBUF_X2 inst_17343 ( .A(net_17190), .Z(net_17191) );
SDFF_X2 inst_1948 ( .D(net_7274), .SI(net_6931), .Q(net_6931), .SE(net_6281), .CK(net_17342) );
DFFR_X2 inst_7158 ( .QN(net_5952), .D(net_2860), .CK(net_16158), .RN(x6501) );
AOI22_X2 inst_8409 ( .B1(net_8860), .A1(net_8305), .B2(net_6252), .A2(net_4345), .ZN(net_3643) );
CLKBUF_X2 inst_15148 ( .A(net_14995), .Z(net_14996) );
AOI22_X2 inst_8266 ( .B1(net_8801), .A1(net_8542), .A2(net_3861), .B2(net_3860), .ZN(net_3772) );
SDFF_X2 inst_422 ( .SI(net_8304), .Q(net_8304), .D(net_3981), .SE(net_3978), .CK(net_13001) );
CLKBUF_X2 inst_16281 ( .A(net_12307), .Z(net_16129) );
SDFFR_X2 inst_2243 ( .SI(net_7388), .SE(net_2814), .Q(net_247), .D(net_247), .CK(net_17454), .RN(x6501) );
SDFF_X2 inst_1426 ( .SI(net_7286), .Q(net_7063), .D(net_7063), .SE(net_6280), .CK(net_16230) );
AOI211_X2 inst_9021 ( .ZN(net_1623), .A(net_1622), .C1(net_1507), .B(net_1503), .C2(net_602) );
NAND2_X2 inst_4812 ( .ZN(net_2912), .A2(net_1282), .A1(net_1266) );
OAI21_X2 inst_3090 ( .B2(net_2897), .ZN(net_2896), .A(net_2844), .B1(net_745) );
CLKBUF_X2 inst_14466 ( .A(net_14313), .Z(net_14314) );
CLKBUF_X2 inst_17050 ( .A(net_16897), .Z(net_16898) );
CLKBUF_X2 inst_14635 ( .A(net_14482), .Z(net_14483) );
CLKBUF_X2 inst_10012 ( .A(net_9859), .Z(net_9860) );
CLKBUF_X2 inst_17751 ( .A(net_17598), .Z(net_17599) );
CLKBUF_X2 inst_14624 ( .A(net_12729), .Z(net_14472) );
AOI22_X2 inst_8355 ( .B1(net_8776), .A1(net_8406), .A2(net_3867), .B2(net_3866), .ZN(net_3693) );
NAND2_X2 inst_4879 ( .ZN(net_791), .A1(net_790), .A2(net_789) );
NAND2_X2 inst_4695 ( .ZN(net_2183), .A2(net_1902), .A1(net_580) );
NAND2_X2 inst_4142 ( .ZN(net_5377), .A1(net_5215), .A2(net_5000) );
CLKBUF_X2 inst_17871 ( .A(net_17718), .Z(net_17719) );
CLKBUF_X2 inst_12125 ( .A(net_11972), .Z(net_11973) );
AOI22_X2 inst_8513 ( .B1(net_6749), .A1(net_6716), .B2(net_6202), .A2(net_3520), .ZN(net_3427) );
CLKBUF_X2 inst_17591 ( .A(net_17438), .Z(net_17439) );
CLKBUF_X2 inst_11260 ( .A(net_11107), .Z(net_11108) );
AND2_X4 inst_9097 ( .ZN(net_2562), .A2(net_2264), .A1(net_1371) );
CLKBUF_X2 inst_12680 ( .A(net_12527), .Z(net_12528) );
CLKBUF_X2 inst_12206 ( .A(net_12053), .Z(net_12054) );
CLKBUF_X2 inst_15267 ( .A(net_15114), .Z(net_15115) );
CLKBUF_X2 inst_14774 ( .A(net_14621), .Z(net_14622) );
OR2_X4 inst_2859 ( .ZN(net_6277), .A1(net_2200), .A2(net_2192) );
CLKBUF_X2 inst_18036 ( .A(net_16270), .Z(net_17884) );
SDFF_X2 inst_397 ( .SI(net_8308), .Q(net_8308), .SE(net_3978), .D(net_3962), .CK(net_10203) );
SDFF_X2 inst_504 ( .SI(net_8597), .Q(net_8597), .SE(net_3984), .D(net_3938), .CK(net_13056) );
AOI222_X1 inst_8601 ( .B2(net_6762), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5823), .A1(net_2149), .C1(x3372) );
CLKBUF_X2 inst_14240 ( .A(net_14087), .Z(net_14088) );
SDFF_X2 inst_1297 ( .SI(net_7672), .Q(net_7672), .SE(net_2714), .D(net_2705), .CK(net_18575) );
OAI211_X2 inst_3194 ( .ZN(net_3219), .C2(net_3161), .B(net_3005), .A(net_2452), .C1(net_1303) );
NAND3_X2 inst_3884 ( .ZN(net_5887), .A3(net_5774), .A1(net_4961), .A2(net_4782) );
CLKBUF_X2 inst_13831 ( .A(net_13678), .Z(net_13679) );
CLKBUF_X2 inst_16937 ( .A(net_9823), .Z(net_16785) );
INV_X2 inst_6296 ( .ZN(net_4202), .A(net_3911) );
SDFF_X2 inst_1173 ( .D(net_7322), .SI(net_6498), .Q(net_6498), .SE(net_3071), .CK(net_9149) );
CLKBUF_X2 inst_9708 ( .A(net_9202), .Z(net_9556) );
OAI22_X2 inst_2908 ( .A2(net_8229), .B2(net_6132), .A1(net_4954), .ZN(net_4876), .B1(net_1395) );
INV_X8 inst_5019 ( .ZN(net_5654), .A(net_4950) );
CLKBUF_X2 inst_9507 ( .A(net_9354), .Z(net_9355) );
CLKBUF_X2 inst_17438 ( .A(net_17285), .Z(net_17286) );
NAND2_X2 inst_4893 ( .A2(net_7525), .A1(net_7522), .ZN(net_1661) );
INV_X4 inst_5875 ( .A(net_7418), .ZN(net_1763) );
CLKBUF_X2 inst_11318 ( .A(net_9712), .Z(net_11166) );
AOI22_X2 inst_8514 ( .B1(net_6683), .A1(net_6650), .A2(net_6213), .B2(net_6138), .ZN(net_3426) );
DFF_X1 inst_6717 ( .QN(net_6794), .D(net_5619), .CK(net_11593) );
CLKBUF_X2 inst_17070 ( .A(net_12211), .Z(net_16918) );
CLKBUF_X2 inst_9807 ( .A(net_9452), .Z(net_9655) );
AND2_X4 inst_9089 ( .A1(net_6120), .ZN(net_4799), .A2(net_2474) );
CLKBUF_X2 inst_13684 ( .A(net_13531), .Z(net_13532) );
CLKBUF_X2 inst_9302 ( .A(net_9145), .Z(net_9150) );
CLKBUF_X2 inst_12995 ( .A(net_12842), .Z(net_12843) );
INV_X2 inst_6283 ( .ZN(net_4218), .A(net_3931) );
DFFR_X1 inst_7380 ( .D(net_5911), .CK(net_17189), .RN(x6501), .Q(x240) );
DFFR_X1 inst_7387 ( .D(net_5846), .CK(net_17179), .RN(x6501), .Q(x291) );
INV_X4 inst_5857 ( .A(net_7562), .ZN(net_3138) );
CLKBUF_X2 inst_9463 ( .A(net_9146), .Z(net_9311) );
SDFF_X2 inst_1774 ( .D(net_7279), .SI(net_6976), .Q(net_6976), .SE(net_6283), .CK(net_14630) );
AOI22_X2 inst_8032 ( .B1(net_8135), .A1(net_7897), .A2(net_6098), .B2(net_4190), .ZN(net_4106) );
CLKBUF_X2 inst_12596 ( .A(net_10853), .Z(net_12444) );
SDFF_X2 inst_985 ( .D(net_7321), .SI(net_6629), .Q(net_6629), .SE(net_3123), .CK(net_12117) );
CLKBUF_X2 inst_12473 ( .A(net_12320), .Z(net_12321) );
DFFS_X1 inst_6943 ( .D(net_6145), .CK(net_13637), .SN(x6501), .Q(x764) );
CLKBUF_X2 inst_16202 ( .A(net_16049), .Z(net_16050) );
CLKBUF_X2 inst_12985 ( .A(net_12832), .Z(net_12833) );
CLKBUF_X2 inst_10627 ( .A(net_10114), .Z(net_10475) );
CLKBUF_X2 inst_17408 ( .A(net_17255), .Z(net_17256) );
CLKBUF_X2 inst_14208 ( .A(net_14055), .Z(net_14056) );
CLKBUF_X2 inst_12563 ( .A(net_12410), .Z(net_12411) );
INV_X4 inst_5918 ( .A(net_6401), .ZN(net_818) );
CLKBUF_X2 inst_12969 ( .A(net_12816), .Z(net_12817) );
SDFF_X2 inst_2007 ( .SI(net_7798), .Q(net_7798), .D(net_2710), .SE(net_2459), .CK(net_14386) );
NAND4_X2 inst_3644 ( .ZN(net_4917), .A3(net_4676), .A2(net_4552), .A4(net_4550), .A1(net_4466) );
CLKBUF_X2 inst_10965 ( .A(net_10812), .Z(net_10813) );
SDFF_X2 inst_805 ( .SI(net_8493), .Q(net_8493), .D(net_3962), .SE(net_3884), .CK(net_10146) );
CLKBUF_X2 inst_9991 ( .A(net_9838), .Z(net_9839) );
INV_X4 inst_6005 ( .A(net_8282), .ZN(net_955) );
CLKBUF_X2 inst_17822 ( .A(net_10106), .Z(net_17670) );
CLKBUF_X2 inst_12387 ( .A(net_12234), .Z(net_12235) );
CLKBUF_X2 inst_12664 ( .A(net_12511), .Z(net_12512) );
CLKBUF_X2 inst_13735 ( .A(net_13582), .Z(net_13583) );
INV_X4 inst_5603 ( .A(net_7386), .ZN(net_643) );
CLKBUF_X2 inst_14257 ( .A(net_14104), .Z(net_14105) );
INV_X2 inst_6569 ( .ZN(net_1653), .A(x5001) );
SDFF_X2 inst_373 ( .SI(net_8313), .Q(net_8313), .SE(net_3978), .D(net_3944), .CK(net_12295) );
CLKBUF_X2 inst_17801 ( .A(net_16300), .Z(net_17649) );
SDFF_X2 inst_1868 ( .D(net_7269), .SI(net_6926), .Q(net_6926), .SE(net_6281), .CK(net_14106) );
CLKBUF_X2 inst_13672 ( .A(net_13421), .Z(net_13520) );
CLKBUF_X2 inst_11428 ( .A(net_10643), .Z(net_11276) );
CLKBUF_X2 inst_9537 ( .A(net_9285), .Z(net_9385) );
XOR2_X2 inst_22 ( .Z(net_1396), .B(net_1395), .A(net_650) );
CLKBUF_X2 inst_19139 ( .A(net_18986), .Z(net_18987) );
CLKBUF_X2 inst_13914 ( .A(net_13761), .Z(net_13762) );
OAI21_X2 inst_3099 ( .ZN(net_2766), .A(net_2765), .B1(net_2764), .B2(net_2048) );
CLKBUF_X2 inst_13289 ( .A(net_9506), .Z(net_13137) );
DFFR_X2 inst_7034 ( .QN(net_7493), .D(net_5039), .CK(net_17256), .RN(x6501) );
SDFF_X2 inst_767 ( .Q(net_8810), .D(net_8810), .SI(net_3950), .SE(net_3879), .CK(net_12588) );
CLKBUF_X2 inst_14065 ( .A(net_9656), .Z(net_13913) );
NOR2_X2 inst_3356 ( .ZN(net_5569), .A2(net_5404), .A1(net_5403) );
CLKBUF_X2 inst_10405 ( .A(net_9512), .Z(net_10253) );
CLKBUF_X2 inst_18270 ( .A(net_18117), .Z(net_18118) );
AOI22_X2 inst_7914 ( .B1(net_8973), .B2(net_5456), .A2(net_4501), .ZN(net_4499), .A1(net_2741) );
CLKBUF_X2 inst_15374 ( .A(net_15221), .Z(net_15222) );
NAND2_X2 inst_4310 ( .A1(net_7055), .A2(net_5162), .ZN(net_5147) );
AOI21_X2 inst_8943 ( .B2(net_5784), .ZN(net_5605), .A(net_5602), .B1(net_2675) );
SDFF_X2 inst_526 ( .Q(net_8854), .D(net_8854), .SI(net_3980), .SE(net_3936), .CK(net_13353) );
SDFF_X2 inst_1178 ( .SI(net_7341), .Q(net_6616), .D(net_6616), .SE(net_3069), .CK(net_11855) );
OAI21_X2 inst_3104 ( .B2(net_8254), .ZN(net_2516), .A(net_2409), .B1(net_1137) );
AND2_X2 inst_9174 ( .A2(net_6188), .ZN(net_2504), .A1(net_2393) );
SDFF_X2 inst_1450 ( .SI(net_7302), .Q(net_7119), .D(net_7119), .SE(net_6278), .CK(net_15898) );
AOI22_X2 inst_8423 ( .B1(net_6596), .A1(net_6563), .A2(net_6257), .B2(net_6110), .ZN(net_3518) );
HA_X1 inst_6689 ( .A(net_3056), .S(net_2927), .CO(net_2926), .B(net_2567) );
INV_X4 inst_5511 ( .A(net_1501), .ZN(net_685) );
OAI21_X2 inst_3123 ( .ZN(net_2284), .A(net_2283), .B2(net_2282), .B1(net_1216) );
CLKBUF_X2 inst_11592 ( .A(net_11439), .Z(net_11440) );
CLKBUF_X2 inst_11149 ( .A(net_9428), .Z(net_10997) );
CLKBUF_X2 inst_10645 ( .A(net_10492), .Z(net_10493) );
CLKBUF_X2 inst_16098 ( .A(net_14192), .Z(net_15946) );
NAND4_X2 inst_3725 ( .ZN(net_4305), .A1(net_4166), .A2(net_4165), .A3(net_4164), .A4(net_4163) );
INV_X4 inst_5400 ( .ZN(net_1283), .A(net_1060) );
SDFF_X2 inst_1592 ( .Q(net_8123), .D(net_8123), .SI(net_2706), .SE(net_2541), .CK(net_18043) );
SDFF_X2 inst_1770 ( .D(net_7290), .SI(net_6867), .Q(net_6867), .SE(net_6282), .CK(net_15342) );
NOR2_X2 inst_3413 ( .ZN(net_3315), .A1(net_3221), .A2(net_3220) );
INV_X4 inst_6095 ( .A(net_7603), .ZN(net_1581) );
NAND2_X2 inst_4483 ( .A2(net_5267), .ZN(net_4495), .A1(net_168) );
CLKBUF_X2 inst_12857 ( .A(net_12323), .Z(net_12705) );
CLKBUF_X2 inst_15617 ( .A(net_11005), .Z(net_15465) );
CLKBUF_X2 inst_11109 ( .A(net_10956), .Z(net_10957) );
CLKBUF_X2 inst_14132 ( .A(net_13979), .Z(net_13980) );
CLKBUF_X2 inst_16776 ( .A(net_16623), .Z(net_16624) );
CLKBUF_X2 inst_18734 ( .A(net_18581), .Z(net_18582) );
SDFF_X2 inst_1419 ( .SI(net_7270), .Q(net_7047), .D(net_7047), .SE(net_6280), .CK(net_16864) );
CLKBUF_X2 inst_14544 ( .A(net_10901), .Z(net_14392) );
SDFFR_X2 inst_2501 ( .Q(net_8979), .D(net_8979), .SI(net_2630), .SE(net_2562), .CK(net_13916), .RN(x6501) );
CLKBUF_X2 inst_18665 ( .A(net_18512), .Z(net_18513) );
CLKBUF_X2 inst_14164 ( .A(net_14011), .Z(net_14012) );
CLKBUF_X2 inst_16233 ( .A(net_16080), .Z(net_16081) );
CLKBUF_X2 inst_18796 ( .A(net_14927), .Z(net_18644) );
CLKBUF_X2 inst_16657 ( .A(net_16504), .Z(net_16505) );
CLKBUF_X2 inst_13314 ( .A(net_13161), .Z(net_13162) );
SDFFR_X2 inst_2378 ( .SE(net_2260), .Q(net_327), .D(net_327), .CK(net_10424), .RN(x6501), .SI(x2805) );
CLKBUF_X2 inst_15942 ( .A(net_15789), .Z(net_15790) );
INV_X2 inst_6302 ( .ZN(net_3989), .A(net_3905) );
CLKBUF_X2 inst_14137 ( .A(net_9897), .Z(net_13985) );
CLKBUF_X2 inst_9996 ( .A(net_9092), .Z(net_9844) );
CLKBUF_X2 inst_14392 ( .A(net_10174), .Z(net_14240) );
CLKBUF_X2 inst_13874 ( .A(net_13721), .Z(net_13722) );
CLKBUF_X2 inst_13164 ( .A(net_12578), .Z(net_13012) );
CLKBUF_X2 inst_16472 ( .A(net_14962), .Z(net_16320) );
CLKBUF_X2 inst_12079 ( .A(net_10060), .Z(net_11927) );
CLKBUF_X2 inst_15237 ( .A(net_9796), .Z(net_15085) );
CLKBUF_X2 inst_10072 ( .A(net_9919), .Z(net_9920) );
CLKBUF_X2 inst_17482 ( .A(net_17329), .Z(net_17330) );
CLKBUF_X2 inst_11153 ( .A(net_11000), .Z(net_11001) );
CLKBUF_X2 inst_16885 ( .A(net_16732), .Z(net_16733) );
CLKBUF_X2 inst_16018 ( .A(net_11096), .Z(net_15866) );
CLKBUF_X2 inst_15569 ( .A(net_12156), .Z(net_15417) );
CLKBUF_X2 inst_12031 ( .A(net_11878), .Z(net_11879) );
CLKBUF_X2 inst_14560 ( .A(net_14407), .Z(net_14408) );
DFF_X1 inst_6740 ( .Q(net_6757), .D(net_5629), .CK(net_10440) );
CLKBUF_X2 inst_10501 ( .A(net_9080), .Z(net_10349) );
CLKBUF_X2 inst_10796 ( .A(net_10643), .Z(net_10644) );
AOI221_X2 inst_8847 ( .B1(net_8569), .C1(net_8458), .C2(net_6263), .B2(net_6262), .ZN(net_6241), .A(net_4263) );
CLKBUF_X2 inst_16616 ( .A(net_16463), .Z(net_16464) );
NAND4_X2 inst_3801 ( .ZN(net_3625), .A1(net_3483), .A2(net_3482), .A3(net_3481), .A4(net_3480) );
NAND2_X2 inst_4177 ( .ZN(net_5329), .A2(net_5192), .A1(net_5078) );
CLKBUF_X2 inst_9350 ( .A(net_9153), .Z(net_9198) );
CLKBUF_X2 inst_17187 ( .A(net_17034), .Z(net_17035) );
INV_X2 inst_6491 ( .A(net_5948), .ZN(net_553) );
CLKBUF_X2 inst_15870 ( .A(net_12050), .Z(net_15718) );
CLKBUF_X2 inst_13133 ( .A(net_12980), .Z(net_12981) );
AND2_X2 inst_9193 ( .ZN(net_1761), .A1(net_1583), .A2(net_1582) );
SDFFR_X2 inst_2155 ( .Q(net_8278), .D(net_8278), .SI(net_8274), .SE(net_2996), .CK(net_18438), .RN(x6501) );
CLKBUF_X2 inst_12927 ( .A(net_12774), .Z(net_12775) );
INV_X2 inst_6352 ( .ZN(net_2257), .A(net_2189) );
SDFF_X2 inst_464 ( .SI(net_8468), .Q(net_8468), .SE(net_3983), .D(net_3942), .CK(net_10081) );
CLKBUF_X2 inst_13428 ( .A(net_13275), .Z(net_13276) );
INV_X4 inst_5360 ( .ZN(net_2803), .A(net_1144) );
CLKBUF_X2 inst_13392 ( .A(net_13239), .Z(net_13240) );
SDFF_X2 inst_341 ( .SI(net_8606), .Q(net_8606), .SE(net_3984), .D(net_3966), .CK(net_10050) );
CLKBUF_X2 inst_15194 ( .A(net_15041), .Z(net_15042) );
CLKBUF_X2 inst_12313 ( .A(net_10154), .Z(net_12161) );
CLKBUF_X2 inst_14961 ( .A(net_13147), .Z(net_14809) );
CLKBUF_X2 inst_13090 ( .A(net_11007), .Z(net_12938) );
CLKBUF_X2 inst_14006 ( .A(net_13853), .Z(net_13854) );
CLKBUF_X2 inst_11095 ( .A(net_9782), .Z(net_10943) );
SDFFR_X2 inst_2359 ( .SE(net_2260), .Q(net_332), .D(net_332), .CK(net_9310), .RN(x6501), .SI(x2542) );
NAND4_X2 inst_3702 ( .ZN(net_4435), .A4(net_4338), .A1(net_3751), .A2(net_3750), .A3(net_3749) );
CLKBUF_X2 inst_11229 ( .A(net_9833), .Z(net_11077) );
AOI22_X2 inst_8526 ( .B1(net_6656), .A1(net_6623), .A2(net_6213), .B2(net_6138), .ZN(net_3414) );
CLKBUF_X2 inst_17090 ( .A(net_16937), .Z(net_16938) );
CLKBUF_X2 inst_13913 ( .A(net_13760), .Z(net_13761) );
CLKBUF_X2 inst_13031 ( .A(net_12878), .Z(net_12879) );
AOI22_X2 inst_8505 ( .B1(net_6720), .A1(net_6687), .B2(net_6202), .A2(net_3520), .ZN(net_3435) );
INV_X4 inst_5556 ( .ZN(net_633), .A(net_632) );
DFF_X1 inst_6826 ( .Q(net_6446), .D(net_3622), .CK(net_17918) );
CLKBUF_X2 inst_10226 ( .A(net_9472), .Z(net_10074) );
CLKBUF_X2 inst_19160 ( .A(net_9300), .Z(net_19008) );
AOI221_X2 inst_8840 ( .C1(net_8150), .B1(net_7708), .C2(net_6101), .B2(net_6095), .ZN(net_6025), .A(net_4282) );
MUX2_X2 inst_4968 ( .S(net_2378), .Z(net_2355), .A(net_1330), .B(net_851) );
CLKBUF_X2 inst_14319 ( .A(net_14166), .Z(net_14167) );
CLKBUF_X2 inst_10122 ( .A(net_9969), .Z(net_9970) );
NAND2_X2 inst_4162 ( .ZN(net_5351), .A2(net_5202), .A1(net_5093) );
INV_X4 inst_5171 ( .A(net_5902), .ZN(net_5824) );
CLKBUF_X2 inst_12936 ( .A(net_10653), .Z(net_12784) );
CLKBUF_X2 inst_18600 ( .A(net_18447), .Z(net_18448) );
CLKBUF_X2 inst_17812 ( .A(net_9234), .Z(net_17660) );
CLKBUF_X2 inst_14363 ( .A(net_12897), .Z(net_14211) );
OAI211_X2 inst_3201 ( .ZN(net_2799), .C2(net_2525), .B(net_2322), .A(net_2202), .C1(net_856) );
CLKBUF_X2 inst_17554 ( .A(net_12992), .Z(net_17402) );
CLKBUF_X2 inst_17930 ( .A(net_17777), .Z(net_17778) );
CLKBUF_X2 inst_14532 ( .A(net_14379), .Z(net_14380) );
CLKBUF_X2 inst_16080 ( .A(net_15927), .Z(net_15928) );
XNOR2_X2 inst_251 ( .B(net_2670), .ZN(net_1199), .A(net_1198) );
CLKBUF_X2 inst_10651 ( .A(net_9335), .Z(net_10499) );
SDFF_X2 inst_1552 ( .Q(net_7979), .D(net_7979), .SI(net_2655), .SE(net_2542), .CK(net_15442) );
SDFF_X2 inst_1524 ( .Q(net_7896), .D(net_7896), .SI(net_2712), .SE(net_2543), .CK(net_17144) );
CLKBUF_X2 inst_18171 ( .A(net_18018), .Z(net_18019) );
CLKBUF_X2 inst_13983 ( .A(net_10996), .Z(net_13831) );
CLKBUF_X2 inst_9369 ( .A(net_9125), .Z(net_9217) );
NAND2_X2 inst_4789 ( .ZN(net_1531), .A2(net_1247), .A1(net_1246) );
MUX2_X2 inst_4977 ( .A(net_9016), .Z(net_3943), .B(net_1468), .S(net_622) );
CLKBUF_X2 inst_15481 ( .A(net_13010), .Z(net_15329) );
CLKBUF_X2 inst_9892 ( .A(net_9187), .Z(net_9740) );
AOI22_X2 inst_7781 ( .A1(net_5268), .ZN(net_4870), .A2(net_4634), .B2(net_4388), .B1(net_2598) );
CLKBUF_X2 inst_18522 ( .A(net_18278), .Z(net_18370) );
CLKBUF_X2 inst_15734 ( .A(net_15581), .Z(net_15582) );
CLKBUF_X2 inst_13628 ( .A(net_13475), .Z(net_13476) );
SDFF_X2 inst_898 ( .SI(net_8714), .Q(net_8714), .SE(net_6195), .D(net_3960), .CK(net_13084) );
SDFF_X2 inst_1977 ( .D(net_7293), .SI(net_6910), .Q(net_6910), .SE(net_6284), .CK(net_18352) );
SDFF_X2 inst_1793 ( .D(net_7283), .SI(net_6980), .Q(net_6980), .SE(net_6283), .CK(net_19015) );
AOI22_X2 inst_8012 ( .B1(net_8098), .A1(net_7758), .B2(net_6108), .A2(net_6096), .ZN(net_4123) );
CLKBUF_X2 inst_9223 ( .A(net_9070), .Z(net_9071) );
CLKBUF_X2 inst_9747 ( .A(net_9594), .Z(net_9595) );
CLKBUF_X2 inst_11804 ( .A(net_11651), .Z(net_11652) );
INV_X4 inst_5299 ( .A(net_1681), .ZN(net_1596) );
CLKBUF_X2 inst_10805 ( .A(net_10652), .Z(net_10653) );
INV_X4 inst_5697 ( .A(net_7365), .ZN(net_1280) );
SDFFR_X2 inst_2291 ( .SE(net_2793), .SI(net_2785), .Q(net_240), .D(net_240), .CK(net_17824), .RN(x6501) );
AOI22_X2 inst_8230 ( .B1(net_8834), .A1(net_8353), .A2(net_6265), .B2(net_6253), .ZN(net_3807) );
NAND2_X2 inst_4822 ( .A1(net_7258), .A2(net_7210), .ZN(net_1520) );
OAI21_X2 inst_3132 ( .ZN(net_2160), .B2(net_2159), .B1(net_2156), .A(net_1351) );
CLKBUF_X2 inst_16572 ( .A(net_13277), .Z(net_16420) );
CLKBUF_X2 inst_13835 ( .A(net_13682), .Z(net_13683) );
CLKBUF_X2 inst_18768 ( .A(net_12621), .Z(net_18616) );
CLKBUF_X2 inst_16419 ( .A(net_16266), .Z(net_16267) );
DFFR_X1 inst_7395 ( .D(net_5834), .CK(net_17175), .RN(x6501), .Q(x275) );
MUX2_X2 inst_4999 ( .A(net_9022), .Z(net_3981), .B(net_747), .S(net_622) );
INV_X4 inst_6071 ( .A(net_6291), .ZN(net_2674) );
INV_X4 inst_5819 ( .A(net_8961), .ZN(net_2039) );
NAND3_X2 inst_3910 ( .ZN(net_5628), .A1(net_5557), .A3(net_5491), .A2(net_5354) );
CLKBUF_X2 inst_18540 ( .A(net_18387), .Z(net_18388) );
SDFF_X2 inst_1332 ( .Q(net_7951), .D(net_7951), .SE(net_2755), .SI(net_2573), .CK(net_18083) );
SDFF_X2 inst_1841 ( .D(net_7292), .SI(net_6909), .Q(net_6909), .SE(net_6284), .CK(net_14886) );
NOR2_X2 inst_3345 ( .ZN(net_5580), .A1(net_5450), .A2(net_5449) );
NOR3_X2 inst_3264 ( .ZN(net_6151), .A1(net_2947), .A2(net_2912), .A3(net_2338) );
CLKBUF_X2 inst_16802 ( .A(net_9537), .Z(net_16650) );
SDFFR_X2 inst_2332 ( .SE(net_2260), .Q(net_353), .D(net_353), .CK(net_9317), .RN(x6501), .SI(x2169) );
CLKBUF_X2 inst_13415 ( .A(net_13262), .Z(net_13263) );
AND2_X4 inst_9082 ( .ZN(net_3069), .A1(net_2904), .A2(net_2903) );
CLKBUF_X2 inst_13431 ( .A(net_13278), .Z(net_13279) );
CLKBUF_X2 inst_18538 ( .A(net_18385), .Z(net_18386) );
CLKBUF_X2 inst_17455 ( .A(net_9360), .Z(net_17303) );
CLKBUF_X2 inst_16019 ( .A(net_13620), .Z(net_15867) );
INV_X4 inst_5946 ( .A(net_8911), .ZN(net_2624) );
SDFFR_X2 inst_2310 ( .SI(net_7407), .SE(net_2260), .Q(net_344), .D(net_344), .CK(net_9366), .RN(x6501) );
CLKBUF_X2 inst_14327 ( .A(net_14174), .Z(net_14175) );
INV_X8 inst_5017 ( .ZN(net_5538), .A(net_4384) );
SDFF_X2 inst_1290 ( .Q(net_8105), .D(net_8105), .SE(net_2707), .SI(net_2639), .CK(net_14437) );
CLKBUF_X2 inst_16461 ( .A(net_11096), .Z(net_16309) );
AOI22_X2 inst_7939 ( .B1(net_8089), .A1(net_7749), .B2(net_6108), .A2(net_6096), .ZN(net_4186) );
CLKBUF_X2 inst_11451 ( .A(net_11298), .Z(net_11299) );
INV_X2 inst_6342 ( .ZN(net_2511), .A(net_2510) );
INV_X4 inst_5845 ( .A(net_7383), .ZN(net_1026) );
INV_X8 inst_5038 ( .ZN(net_6095), .A(net_3576) );
CLKBUF_X2 inst_18090 ( .A(net_17937), .Z(net_17938) );
CLKBUF_X2 inst_13399 ( .A(net_13246), .Z(net_13247) );
INV_X4 inst_5142 ( .A(net_3888), .ZN(net_3599) );
INV_X4 inst_5757 ( .A(net_8889), .ZN(net_3587) );
NAND2_X2 inst_4899 ( .A2(net_7394), .ZN(net_621), .A1(net_183) );
CLKBUF_X2 inst_15865 ( .A(net_15712), .Z(net_15713) );
CLKBUF_X2 inst_12604 ( .A(net_12451), .Z(net_12452) );
INV_X4 inst_5079 ( .ZN(net_5842), .A(net_5789) );
INV_X2 inst_6429 ( .ZN(net_715), .A(net_714) );
NAND4_X2 inst_3861 ( .A2(net_4465), .A3(net_4459), .A1(net_4457), .A4(net_3236), .ZN(net_1442) );
CLKBUF_X2 inst_15809 ( .A(net_15656), .Z(net_15657) );
NAND2_X2 inst_4399 ( .A1(net_7086), .A2(net_5164), .ZN(net_5058) );
CLKBUF_X2 inst_11547 ( .A(net_11394), .Z(net_11395) );
CLKBUF_X2 inst_9847 ( .A(net_9694), .Z(net_9695) );
CLKBUF_X2 inst_9840 ( .A(net_9258), .Z(net_9688) );
CLKBUF_X2 inst_16864 ( .A(net_16711), .Z(net_16712) );
NAND2_X2 inst_4196 ( .ZN(net_5302), .A1(net_5179), .A2(net_4982) );
CLKBUF_X2 inst_10672 ( .A(net_10519), .Z(net_10520) );
SDFF_X2 inst_1014 ( .SI(net_7328), .Q(net_6669), .D(net_6669), .SE(net_3126), .CK(net_9520) );
SDFFR_X2 inst_2531 ( .Q(net_7668), .D(net_7668), .SE(net_2299), .SI(net_1579), .CK(net_17439), .RN(x6501) );
CLKBUF_X2 inst_10009 ( .A(net_9856), .Z(net_9857) );
DFF_X1 inst_6781 ( .Q(net_7530), .D(net_4589), .CK(net_9394) );
CLKBUF_X2 inst_14918 ( .A(net_14765), .Z(net_14766) );
CLKBUF_X2 inst_11879 ( .A(net_11726), .Z(net_11727) );
CLKBUF_X2 inst_16597 ( .A(net_16444), .Z(net_16445) );
CLKBUF_X2 inst_18363 ( .A(net_12957), .Z(net_18211) );
CLKBUF_X2 inst_12299 ( .A(net_10796), .Z(net_12147) );
CLKBUF_X2 inst_16479 ( .A(net_11254), .Z(net_16327) );
SDFF_X2 inst_1680 ( .Q(net_8149), .D(net_8149), .SI(net_2655), .SE(net_2538), .CK(net_15496) );
CLKBUF_X2 inst_15221 ( .A(net_11409), .Z(net_15069) );
SDFF_X2 inst_1626 ( .Q(net_8170), .D(net_8170), .SI(net_2717), .SE(net_2538), .CK(net_16479) );
CLKBUF_X2 inst_12834 ( .A(net_11271), .Z(net_12682) );
CLKBUF_X2 inst_16323 ( .A(net_16170), .Z(net_16171) );
CLKBUF_X2 inst_12271 ( .A(net_12118), .Z(net_12119) );
INV_X2 inst_6528 ( .A(net_6377), .ZN(net_2144) );
CLKBUF_X2 inst_9789 ( .A(net_9636), .Z(net_9637) );
AND2_X4 inst_9117 ( .A1(net_7405), .ZN(net_1703), .A2(net_1347) );
NAND3_X2 inst_3894 ( .ZN(net_5644), .A1(net_5573), .A3(net_5507), .A2(net_5418) );
AOI22_X2 inst_8037 ( .A1(net_7966), .B1(net_7796), .A2(net_6092), .B2(net_6091), .ZN(net_4102) );
CLKBUF_X2 inst_10132 ( .A(net_9979), .Z(net_9980) );
INV_X4 inst_5385 ( .A(net_1149), .ZN(net_1100) );
SDFF_X2 inst_1087 ( .D(net_7341), .SI(net_6517), .Q(net_6517), .SE(net_3071), .CK(net_11879) );
CLKBUF_X2 inst_17055 ( .A(net_10364), .Z(net_16903) );
CLKBUF_X2 inst_13701 ( .A(net_13548), .Z(net_13549) );
CLKBUF_X2 inst_14453 ( .A(net_14300), .Z(net_14301) );
CLKBUF_X2 inst_10061 ( .A(net_9908), .Z(net_9909) );
SDFF_X2 inst_1375 ( .SI(net_7708), .Q(net_7708), .D(net_2709), .SE(net_2559), .CK(net_15774) );
CLKBUF_X2 inst_12199 ( .A(net_9744), .Z(net_12047) );
CLKBUF_X2 inst_15693 ( .A(net_9185), .Z(net_15541) );
AOI22_X2 inst_7966 ( .B1(net_8059), .A1(net_7855), .B2(net_6107), .ZN(net_6004), .A2(net_4400) );
CLKBUF_X2 inst_19097 ( .A(net_18944), .Z(net_18945) );
NAND2_X2 inst_4564 ( .A2(net_7653), .A1(net_6175), .ZN(net_6081) );
CLKBUF_X2 inst_15134 ( .A(net_14981), .Z(net_14982) );
CLKBUF_X2 inst_9290 ( .A(net_9132), .Z(net_9138) );
INV_X4 inst_5258 ( .A(net_2068), .ZN(net_1777) );
CLKBUF_X2 inst_12235 ( .A(net_11640), .Z(net_12083) );
CLKBUF_X2 inst_11209 ( .A(net_11056), .Z(net_11057) );
SDFFR_X2 inst_2564 ( .QN(net_6365), .SE(net_2147), .SI(net_1961), .D(net_697), .CK(net_18130), .RN(x6501) );
CLKBUF_X2 inst_15173 ( .A(net_10048), .Z(net_15021) );
SDFF_X2 inst_1082 ( .D(net_7334), .SI(net_6510), .Q(net_6510), .SE(net_3071), .CK(net_9757) );
CLKBUF_X2 inst_15185 ( .A(net_12087), .Z(net_15033) );
SDFFR_X1 inst_2677 ( .SI(net_7542), .SE(net_5043), .CK(net_9708), .RN(x6501), .Q(x4036), .D(x4036) );
CLKBUF_X2 inst_10068 ( .A(net_9915), .Z(net_9916) );
XOR2_X1 inst_105 ( .A(net_7579), .B(net_3098), .Z(net_995) );
CLKBUF_X2 inst_18529 ( .A(net_18376), .Z(net_18377) );
NOR2_X2 inst_3518 ( .ZN(net_1933), .A1(net_1756), .A2(net_1755) );
CLKBUF_X2 inst_18888 ( .A(net_18735), .Z(net_18736) );
SDFFR_X2 inst_2161 ( .QN(net_7578), .D(net_3967), .SE(net_3144), .SI(net_3140), .CK(net_10876), .RN(x6501) );
AOI22_X2 inst_8294 ( .B1(net_8805), .A1(net_8546), .A2(net_3861), .B2(net_3860), .ZN(net_3748) );
SDFF_X2 inst_625 ( .SI(net_8537), .Q(net_8537), .SE(net_3979), .D(net_3958), .CK(net_13191) );
CLKBUF_X2 inst_16855 ( .A(net_11793), .Z(net_16703) );
DFF_X1 inst_6747 ( .QN(net_6792), .D(net_5621), .CK(net_9545) );
CLKBUF_X2 inst_14041 ( .A(net_13888), .Z(net_13889) );
AOI22_X2 inst_8119 ( .B1(net_8048), .A1(net_7844), .B2(net_6107), .ZN(net_6026), .A2(net_4400) );
XNOR2_X2 inst_181 ( .B(net_5974), .ZN(net_1675), .A(net_1332) );
CLKBUF_X2 inst_17460 ( .A(net_15960), .Z(net_17308) );
CLKBUF_X2 inst_13212 ( .A(net_13059), .Z(net_13060) );
AOI21_X2 inst_8964 ( .ZN(net_3183), .A(net_3182), .B2(net_3181), .B1(x933) );
AOI22_X2 inst_8329 ( .B1(net_8809), .A1(net_8550), .A2(net_3861), .B2(net_3860), .ZN(net_3717) );
INV_X4 inst_5215 ( .ZN(net_2325), .A(net_2324) );
CLKBUF_X2 inst_17470 ( .A(net_9542), .Z(net_17318) );
CLKBUF_X2 inst_17479 ( .A(net_16868), .Z(net_17327) );
CLKBUF_X2 inst_10885 ( .A(net_10732), .Z(net_10733) );
CLKBUF_X2 inst_16723 ( .A(net_16570), .Z(net_16571) );
CLKBUF_X2 inst_18568 ( .A(net_16807), .Z(net_18416) );
CLKBUF_X2 inst_9738 ( .A(net_9585), .Z(net_9586) );
SDFF_X2 inst_713 ( .SI(net_8662), .Q(net_8662), .D(net_3950), .SE(net_3885), .CK(net_10996) );
CLKBUF_X2 inst_10125 ( .A(net_9972), .Z(net_9973) );
CLKBUF_X2 inst_16548 ( .A(net_10103), .Z(net_16396) );
DFFS_X1 inst_6918 ( .D(net_4402), .CK(net_13811), .SN(x6501), .Q(x34) );
CLKBUF_X2 inst_19176 ( .A(net_19023), .Z(net_19024) );
CLKBUF_X2 inst_17578 ( .A(net_15458), .Z(net_17426) );
CLKBUF_X2 inst_11508 ( .A(net_11355), .Z(net_11356) );
CLKBUF_X2 inst_16492 ( .A(net_16339), .Z(net_16340) );
CLKBUF_X2 inst_15256 ( .A(net_15103), .Z(net_15104) );
AOI22_X2 inst_7768 ( .B1(net_6995), .A1(net_6955), .A2(net_5443), .B2(net_5442), .ZN(net_5333) );
CLKBUF_X2 inst_17036 ( .A(net_16883), .Z(net_16884) );
CLKBUF_X2 inst_14062 ( .A(net_13909), .Z(net_13910) );
OAI211_X2 inst_3208 ( .ZN(net_2522), .C1(net_2205), .C2(net_2204), .B(net_2102), .A(net_1754) );
DFFR_X1 inst_7410 ( .D(net_5703), .CK(net_17163), .RN(x6501), .Q(x324) );
NAND2_X2 inst_4134 ( .ZN(net_5388), .A2(net_5220), .A1(net_5120) );
NOR2_X2 inst_3507 ( .A2(net_2400), .ZN(net_2116), .A1(net_1461) );
XNOR2_X2 inst_271 ( .B(net_1444), .ZN(net_1047), .A(net_503) );
CLKBUF_X2 inst_11918 ( .A(net_11710), .Z(net_11766) );
HA_X1 inst_6705 ( .A(net_8261), .S(net_1697), .CO(net_1696), .B(net_1230) );
SDFF_X2 inst_1230 ( .Q(net_7819), .D(net_7819), .SE(net_2730), .SI(net_2720), .CK(net_18096) );
CLKBUF_X2 inst_16979 ( .A(net_16826), .Z(net_16827) );
CLKBUF_X2 inst_10844 ( .A(net_10691), .Z(net_10692) );
DFFR_X2 inst_7262 ( .QN(net_7229), .D(net_1986), .CK(net_14781), .RN(x6501) );
NOR2_X2 inst_3535 ( .ZN(net_1752), .A1(net_1575), .A2(net_1574) );
CLKBUF_X2 inst_17880 ( .A(net_17727), .Z(net_17728) );
CLKBUF_X2 inst_9344 ( .A(net_9191), .Z(net_9192) );
CLKBUF_X2 inst_14685 ( .A(net_14325), .Z(net_14533) );
NOR2_X2 inst_3497 ( .A2(net_2767), .ZN(net_1990), .A1(net_1131) );
CLKBUF_X2 inst_17752 ( .A(net_17599), .Z(net_17600) );
SDFF_X2 inst_1064 ( .D(net_7325), .SI(net_6534), .Q(net_6534), .SE(net_3086), .CK(net_9128) );
INV_X4 inst_5416 ( .ZN(net_3363), .A(net_1075) );
CLKBUF_X2 inst_17193 ( .A(net_12129), .Z(net_17041) );
CLKBUF_X2 inst_14875 ( .A(net_14722), .Z(net_14723) );
CLKBUF_X2 inst_11110 ( .A(net_10957), .Z(net_10958) );
NOR2_X2 inst_3599 ( .ZN(net_1173), .A2(net_845), .A1(net_543) );
CLKBUF_X2 inst_14335 ( .A(net_12558), .Z(net_14183) );
CLKBUF_X2 inst_14539 ( .A(net_10795), .Z(net_14387) );
CLKBUF_X2 inst_17490 ( .A(net_17337), .Z(net_17338) );
CLKBUF_X2 inst_13727 ( .A(net_9157), .Z(net_13575) );
CLKBUF_X2 inst_17737 ( .A(net_14284), .Z(net_17585) );
CLKBUF_X2 inst_12124 ( .A(net_10368), .Z(net_11972) );
INV_X4 inst_5208 ( .A(net_2464), .ZN(net_2383) );
NOR2_X2 inst_3581 ( .A1(net_8217), .ZN(net_2263), .A2(net_759) );
CLKBUF_X2 inst_9930 ( .A(net_9777), .Z(net_9778) );
NAND2_X2 inst_4833 ( .ZN(net_1669), .A2(net_1062), .A1(x12843) );
SDFFS_X2 inst_2065 ( .SI(net_7394), .SE(net_2417), .Q(net_183), .D(net_183), .CK(net_17502), .SN(x6501) );
CLKBUF_X2 inst_10765 ( .A(net_10612), .Z(net_10613) );
SDFFR_X2 inst_2251 ( .D(net_2803), .SE(net_2797), .SI(net_195), .Q(net_195), .CK(net_14986), .RN(x6501) );
NAND3_X2 inst_3987 ( .ZN(net_1735), .A2(net_1422), .A1(net_1398), .A3(net_1384) );
CLKBUF_X2 inst_18008 ( .A(net_9586), .Z(net_17856) );
CLKBUF_X2 inst_12825 ( .A(net_9182), .Z(net_12673) );
CLKBUF_X2 inst_13720 ( .A(net_13567), .Z(net_13568) );
INV_X4 inst_5124 ( .ZN(net_4647), .A(net_4414) );
CLKBUF_X2 inst_18797 ( .A(net_18644), .Z(net_18645) );
CLKBUF_X2 inst_13226 ( .A(net_10898), .Z(net_13074) );
SDFF_X2 inst_1899 ( .D(net_7291), .SI(net_7028), .Q(net_7028), .SE(net_6277), .CK(net_15314) );
DFFR_X2 inst_7200 ( .D(net_2371), .QN(net_218), .CK(net_17568), .RN(x6501) );
CLKBUF_X2 inst_9349 ( .A(net_9196), .Z(net_9197) );
SDFFR_X2 inst_2569 ( .QN(net_6356), .SE(net_2147), .D(net_2121), .SI(net_1808), .CK(net_17523), .RN(x6501) );
CLKBUF_X2 inst_10573 ( .A(net_9972), .Z(net_10421) );
CLKBUF_X2 inst_10197 ( .A(net_10044), .Z(net_10045) );
AND3_X2 inst_9048 ( .A1(net_2346), .ZN(net_1865), .A2(net_1861), .A3(net_1704) );
CLKBUF_X2 inst_19113 ( .A(net_18960), .Z(net_18961) );
SDFFR_X1 inst_2716 ( .SI(net_9015), .Q(net_9015), .D(net_7444), .SE(net_3208), .CK(net_10110), .RN(x6501) );
CLKBUF_X2 inst_17529 ( .A(net_15122), .Z(net_17377) );
NOR4_X2 inst_3228 ( .ZN(net_2276), .A4(net_2004), .A3(net_1967), .A2(net_1015), .A1(net_968) );
CLKBUF_X2 inst_9212 ( .A(net_9059), .Z(net_9060) );
SDFFR_X2 inst_2124 ( .SI(net_7188), .Q(net_7188), .D(net_6439), .SE(net_4362), .CK(net_17840), .RN(x6501) );
CLKBUF_X2 inst_13268 ( .A(net_13115), .Z(net_13116) );
CLKBUF_X2 inst_17095 ( .A(net_16942), .Z(net_16943) );
SDFF_X2 inst_1435 ( .SI(net_7276), .Q(net_7093), .D(net_7093), .SE(net_6278), .CK(net_14141) );
CLKBUF_X2 inst_11582 ( .A(net_11429), .Z(net_11430) );
NAND4_X2 inst_3746 ( .ZN(net_4284), .A1(net_4039), .A2(net_4038), .A3(net_4037), .A4(net_4036) );
CLKBUF_X2 inst_15610 ( .A(net_12441), .Z(net_15458) );
CLKBUF_X2 inst_12288 ( .A(net_12135), .Z(net_12136) );
CLKBUF_X2 inst_10810 ( .A(net_10577), .Z(net_10658) );
NAND2_X2 inst_4121 ( .ZN(net_5405), .A1(net_5229), .A2(net_5007) );
SDFFR_X2 inst_2640 ( .Q(net_7389), .D(net_7389), .SE(net_1136), .CK(net_15863), .RN(x6501), .SI(x4561) );
CLKBUF_X2 inst_16588 ( .A(net_16435), .Z(net_16436) );
CLKBUF_X2 inst_12732 ( .A(net_10212), .Z(net_12580) );
AOI22_X2 inst_8162 ( .B1(net_8667), .A1(net_8630), .B2(net_6109), .ZN(net_3872), .A2(net_3857) );
CLKBUF_X2 inst_18184 ( .A(net_18031), .Z(net_18032) );
AOI22_X2 inst_7908 ( .B1(net_7194), .A2(net_6445), .B2(net_5655), .A1(net_5654), .ZN(net_4517) );
NAND2_X2 inst_4448 ( .A1(net_6848), .A2(net_5016), .ZN(net_4979) );
CLKBUF_X2 inst_17042 ( .A(net_16889), .Z(net_16890) );
CLKBUF_X2 inst_17642 ( .A(net_11234), .Z(net_17490) );
CLKBUF_X2 inst_18941 ( .A(net_18788), .Z(net_18789) );
NAND2_X2 inst_4784 ( .ZN(net_1537), .A1(net_1536), .A2(net_1277) );
CLKBUF_X2 inst_17998 ( .A(net_14536), .Z(net_17846) );
CLKBUF_X2 inst_15155 ( .A(net_15002), .Z(net_15003) );
DFFR_X2 inst_7207 ( .D(net_2365), .QN(net_209), .CK(net_15006), .RN(x6501) );
CLKBUF_X2 inst_12256 ( .A(net_12103), .Z(net_12104) );
CLKBUF_X2 inst_14716 ( .A(net_14563), .Z(net_14564) );
NOR3_X2 inst_3321 ( .A3(net_6406), .ZN(net_2991), .A1(net_1843), .A2(net_1076) );
CLKBUF_X2 inst_16464 ( .A(net_16311), .Z(net_16312) );
XNOR2_X2 inst_333 ( .B(net_7638), .A(net_7635), .ZN(net_794) );
INV_X4 inst_5988 ( .A(net_7438), .ZN(net_3224) );
AOI22_X2 inst_8368 ( .B1(net_8707), .A1(net_8485), .B2(net_4350), .A2(net_4349), .ZN(net_3680) );
CLKBUF_X2 inst_18069 ( .A(net_17916), .Z(net_17917) );
INV_X4 inst_5279 ( .A(net_2397), .ZN(net_1771) );
CLKBUF_X2 inst_11934 ( .A(net_11781), .Z(net_11782) );
CLKBUF_X2 inst_11394 ( .A(net_11241), .Z(net_11242) );
CLKBUF_X2 inst_9335 ( .A(net_9182), .Z(net_9183) );
CLKBUF_X2 inst_10953 ( .A(net_9834), .Z(net_10801) );
CLKBUF_X2 inst_10897 ( .A(net_9123), .Z(net_10745) );
SDFFR_X1 inst_2764 ( .QN(net_7584), .D(net_3942), .SE(net_3144), .SI(net_3107), .CK(net_12661), .RN(x6501) );
INV_X2 inst_6246 ( .ZN(net_4860), .A(net_4754) );
CLKBUF_X2 inst_13755 ( .A(net_9600), .Z(net_13603) );
CLKBUF_X2 inst_17722 ( .A(net_17569), .Z(net_17570) );
CLKBUF_X2 inst_11065 ( .A(net_10912), .Z(net_10913) );
INV_X4 inst_6155 ( .ZN(net_6189), .A(net_4416) );
INV_X4 inst_5774 ( .A(net_7598), .ZN(net_555) );
CLKBUF_X2 inst_9664 ( .A(net_9315), .Z(net_9512) );
AOI221_X4 inst_8719 ( .B1(net_8719), .C1(net_8497), .B2(net_4350), .C2(net_4349), .ZN(net_4348), .A(net_4261) );
CLKBUF_X2 inst_11610 ( .A(net_9545), .Z(net_11458) );
OAI211_X2 inst_3178 ( .ZN(net_5782), .B(net_5747), .C2(net_5534), .C1(net_5452), .A(net_2963) );
NAND2_X2 inst_4203 ( .ZN(net_5293), .A1(net_5053), .A2(net_5052) );
CLKBUF_X2 inst_9972 ( .A(net_9505), .Z(net_9820) );
OR2_X4 inst_2840 ( .A2(net_2290), .ZN(net_2212), .A1(net_2112) );
CLKBUF_X2 inst_16313 ( .A(net_16160), .Z(net_16161) );
CLKBUF_X2 inst_12521 ( .A(net_12368), .Z(net_12369) );
CLKBUF_X2 inst_10939 ( .A(net_10786), .Z(net_10787) );
CLKBUF_X2 inst_14214 ( .A(net_14061), .Z(net_14062) );
SDFFR_X1 inst_2781 ( .D(net_7384), .Q(net_7281), .SI(net_1942), .SE(net_1327), .CK(net_14772), .RN(x6501) );
CLKBUF_X2 inst_9544 ( .A(net_9391), .Z(net_9392) );
CLKBUF_X2 inst_13190 ( .A(net_13037), .Z(net_13038) );
CLKBUF_X2 inst_11043 ( .A(net_10890), .Z(net_10891) );
CLKBUF_X2 inst_18262 ( .A(net_18109), .Z(net_18110) );
CLKBUF_X2 inst_12780 ( .A(net_12439), .Z(net_12628) );
SDFFR_X2 inst_2402 ( .SI(net_7372), .SE(net_2732), .D(net_2695), .QN(net_147), .CK(net_16104), .RN(x6501) );
CLKBUF_X2 inst_18245 ( .A(net_18092), .Z(net_18093) );
AOI21_X2 inst_8877 ( .B2(net_5871), .ZN(net_5868), .A(net_5863), .B1(net_2676) );
SDFFR_X2 inst_2616 ( .Q(net_7368), .D(net_7368), .SE(net_1136), .CK(net_18636), .RN(x6501), .SI(x4840) );
CLKBUF_X2 inst_17701 ( .A(net_17548), .Z(net_17549) );
CLKBUF_X2 inst_14627 ( .A(net_14474), .Z(net_14475) );
AOI22_X2 inst_8095 ( .B1(net_8075), .A1(net_7871), .B2(net_6107), .A2(net_4400), .ZN(net_4052) );
SDFFR_X2 inst_2113 ( .QN(net_8907), .SE(net_6144), .D(net_5034), .SI(net_5033), .CK(net_17586), .RN(x6501) );
INV_X4 inst_5249 ( .ZN(net_2159), .A(net_1769) );
SDFF_X2 inst_1820 ( .D(net_7265), .SI(net_6922), .Q(net_6922), .SE(net_6281), .CK(net_14352) );
CLKBUF_X2 inst_15674 ( .A(net_12845), .Z(net_15522) );
AOI22_X2 inst_8253 ( .B1(net_8762), .A1(net_8392), .A2(net_3867), .B2(net_3866), .ZN(net_3784) );
DFFR_X2 inst_6998 ( .QN(net_5968), .D(net_5875), .CK(net_11546), .RN(x6501) );
INV_X4 inst_6065 ( .A(net_8284), .ZN(net_1020) );
NAND2_X2 inst_4729 ( .ZN(net_2655), .A2(net_1586), .A1(net_1007) );
SDFFR_X2 inst_2271 ( .SI(net_7382), .SE(net_2814), .Q(net_241), .D(net_241), .CK(net_17769), .RN(x6501) );
INV_X2 inst_6209 ( .ZN(net_5501), .A(net_5393) );
AOI22_X2 inst_7793 ( .A2(net_6187), .B2(net_5463), .ZN(net_4805), .B1(net_442), .A1(net_205) );
CLKBUF_X2 inst_16119 ( .A(net_15966), .Z(net_15967) );
CLKBUF_X2 inst_10314 ( .A(net_9489), .Z(net_10162) );
NAND4_X2 inst_3779 ( .ZN(net_4242), .A1(net_3711), .A2(net_3710), .A3(net_3709), .A4(net_3708) );
CLKBUF_X2 inst_11644 ( .A(net_11491), .Z(net_11492) );
SDFF_X2 inst_697 ( .Q(net_8416), .D(net_8416), .SI(net_3937), .SE(net_3934), .CK(net_13035) );
CLKBUF_X2 inst_11150 ( .A(net_10997), .Z(net_10998) );
CLKBUF_X2 inst_14035 ( .A(net_13882), .Z(net_13883) );
INV_X4 inst_5159 ( .ZN(net_6080), .A(net_3180) );
CLKBUF_X2 inst_10350 ( .A(net_10197), .Z(net_10198) );
CLKBUF_X2 inst_18756 ( .A(net_18603), .Z(net_18604) );
DFFR_X1 inst_7527 ( .Q(net_7658), .D(net_7654), .CK(net_12719), .RN(x6501) );
CLKBUF_X2 inst_13941 ( .A(net_13788), .Z(net_13789) );
CLKBUF_X2 inst_11512 ( .A(net_11359), .Z(net_11360) );
CLKBUF_X2 inst_12307 ( .A(net_12154), .Z(net_12155) );
AOI221_X2 inst_8758 ( .C2(net_5609), .B2(net_5520), .ZN(net_5518), .A(net_5026), .C1(net_354), .B1(net_284) );
CLKBUF_X2 inst_12975 ( .A(net_12822), .Z(net_12823) );
CLKBUF_X2 inst_17252 ( .A(net_17099), .Z(net_17100) );
CLKBUF_X2 inst_14853 ( .A(net_14700), .Z(net_14701) );
CLKBUF_X2 inst_13972 ( .A(net_13819), .Z(net_13820) );
CLKBUF_X2 inst_16279 ( .A(net_16126), .Z(net_16127) );
CLKBUF_X2 inst_15165 ( .A(net_15012), .Z(net_15013) );
CLKBUF_X2 inst_14198 ( .A(net_14045), .Z(net_14046) );
CLKBUF_X2 inst_16656 ( .A(net_16503), .Z(net_16504) );
SDFF_X2 inst_2004 ( .SI(net_7787), .Q(net_7787), .D(net_2576), .SE(net_2459), .CK(net_15949) );
CLKBUF_X2 inst_15894 ( .A(net_15644), .Z(net_15742) );
XNOR2_X2 inst_220 ( .ZN(net_1402), .B(net_1401), .A(net_773) );
XNOR2_X2 inst_245 ( .A(net_7571), .B(net_2818), .ZN(net_1213) );
DFFR_X2 inst_6991 ( .QN(net_5972), .D(net_5891), .CK(net_11549), .RN(x6501) );
CLKBUF_X2 inst_9779 ( .A(net_9626), .Z(net_9627) );
CLKBUF_X2 inst_15584 ( .A(net_15431), .Z(net_15432) );
NAND2_X2 inst_4111 ( .ZN(net_5419), .A2(net_5236), .A1(net_5144) );
CLKBUF_X2 inst_19146 ( .A(net_18993), .Z(net_18994) );
AOI22_X2 inst_8388 ( .B1(net_8857), .A1(net_8302), .B2(net_6252), .A2(net_4345), .ZN(net_3660) );
CLKBUF_X2 inst_18164 ( .A(net_17469), .Z(net_18012) );
CLKBUF_X2 inst_16867 ( .A(net_16714), .Z(net_16715) );
AOI221_X2 inst_8768 ( .C1(net_8983), .B2(net_5538), .C2(net_5456), .ZN(net_5280), .A(net_4876), .B1(net_412) );
XNOR2_X2 inst_147 ( .B(net_4714), .ZN(net_2142), .A(net_2037) );
XNOR2_X2 inst_313 ( .B(net_7385), .ZN(net_953), .A(net_558) );
SDFF_X2 inst_1676 ( .SI(net_7746), .Q(net_7746), .D(net_2702), .SE(net_2560), .CK(net_18847) );
NAND2_X2 inst_4170 ( .ZN(net_5340), .A1(net_5086), .A2(net_5085) );
AOI22_X2 inst_8480 ( .B1(net_6543), .A1(net_6510), .A2(net_6137), .B2(net_6104), .ZN(net_3460) );
SDFF_X2 inst_1041 ( .SI(net_7331), .Q(net_6705), .D(net_6705), .SE(net_3125), .CK(net_11291) );
SDFFS_X2 inst_2086 ( .SI(net_7483), .Q(net_7483), .D(net_2760), .SE(net_2340), .CK(net_16092), .SN(x6501) );
CLKBUF_X2 inst_17964 ( .A(net_17811), .Z(net_17812) );
CLKBUF_X2 inst_12918 ( .A(net_12765), .Z(net_12766) );
AOI221_X2 inst_8743 ( .C2(net_6433), .ZN(net_5661), .C1(net_5654), .B2(net_5595), .A(net_5586), .B1(net_315) );
AOI22_X2 inst_8570 ( .A2(net_8251), .A1(net_4729), .B2(net_4728), .B1(net_2786), .ZN(net_2154) );
AOI22_X2 inst_8195 ( .B1(net_8681), .A1(net_8644), .ZN(net_6246), .B2(net_6109), .A2(net_3857) );
CLKBUF_X2 inst_12789 ( .A(net_12636), .Z(net_12637) );
SDFF_X2 inst_553 ( .Q(net_8700), .D(net_8700), .SI(net_3976), .SE(net_3935), .CK(net_12796) );
CLKBUF_X2 inst_9271 ( .A(net_9118), .Z(net_9119) );
NOR2_X4 inst_3331 ( .A2(net_7345), .A1(net_6186), .ZN(net_5984) );
XNOR2_X2 inst_242 ( .B(net_5976), .ZN(net_1219), .A(x3561) );
AOI21_X2 inst_8950 ( .A(net_5783), .ZN(net_5668), .B1(net_5471), .B2(net_5265) );
CLKBUF_X2 inst_16843 ( .A(net_16690), .Z(net_16691) );
CLKBUF_X2 inst_16177 ( .A(net_12986), .Z(net_16025) );
CLKBUF_X2 inst_14592 ( .A(net_14439), .Z(net_14440) );
CLKBUF_X2 inst_16263 ( .A(net_15205), .Z(net_16111) );
SDFF_X2 inst_1186 ( .D(net_7320), .SI(net_6562), .Q(net_6562), .SE(net_3070), .CK(net_9827) );
CLKBUF_X2 inst_9513 ( .A(net_9138), .Z(net_9361) );
CLKBUF_X2 inst_10542 ( .A(net_10389), .Z(net_10390) );
SDFF_X2 inst_1739 ( .SI(net_7269), .Q(net_7126), .D(net_7126), .SE(net_6279), .CK(net_16820) );
CLKBUF_X2 inst_13712 ( .A(net_13559), .Z(net_13560) );
CLKBUF_X2 inst_14863 ( .A(net_14710), .Z(net_14711) );
CLKBUF_X2 inst_12430 ( .A(net_11128), .Z(net_12278) );
INV_X4 inst_5446 ( .A(net_6753), .ZN(net_1465) );
MUX2_X2 inst_4956 ( .A(net_2803), .S(net_2370), .Z(net_2367), .B(net_814) );
NOR2_X2 inst_3609 ( .A2(net_1846), .A1(net_1575), .ZN(net_1169) );
CLKBUF_X2 inst_17631 ( .A(net_17478), .Z(net_17479) );
AOI222_X1 inst_8619 ( .A2(net_8223), .A1(net_4891), .B2(net_4889), .C2(net_4888), .ZN(net_4887), .B1(net_4697), .C1(net_3132) );
CLKBUF_X2 inst_19101 ( .A(net_18948), .Z(net_18949) );
INV_X16 inst_6649 ( .ZN(net_6191), .A(net_6190) );
CLKBUF_X2 inst_13338 ( .A(net_13185), .Z(net_13186) );
CLKBUF_X2 inst_19189 ( .A(net_19036), .Z(net_19037) );
CLKBUF_X2 inst_16809 ( .A(net_16656), .Z(net_16657) );
AOI22_X2 inst_8221 ( .B1(net_8684), .A1(net_8647), .B2(net_6109), .A2(net_3857), .ZN(net_3815) );
SDFFR_X2 inst_2608 ( .D(net_7369), .Q(net_7266), .SI(net_1806), .SE(net_1327), .CK(net_14673), .RN(x6501) );
INV_X4 inst_6008 ( .A(net_8292), .ZN(net_1021) );
CLKBUF_X2 inst_11840 ( .A(net_11687), .Z(net_11688) );
CLKBUF_X2 inst_12659 ( .A(net_12506), .Z(net_12507) );
CLKBUF_X2 inst_15873 ( .A(net_15720), .Z(net_15721) );
CLKBUF_X2 inst_14766 ( .A(net_11119), .Z(net_14614) );
SDFFR_X2 inst_2521 ( .D(net_7369), .SE(net_2387), .SI(net_284), .Q(net_284), .CK(net_16397), .RN(x6501) );
SDFF_X2 inst_385 ( .Q(net_8820), .D(net_8820), .SI(net_3965), .SE(net_3964), .CK(net_13155) );
CLKBUF_X2 inst_14110 ( .A(net_11849), .Z(net_13958) );
SDFFR_X1 inst_2653 ( .D(net_6775), .SE(net_4506), .CK(net_9193), .RN(x6501), .SI(x1639), .Q(x1639) );
CLKBUF_X2 inst_11062 ( .A(net_9502), .Z(net_10910) );
CLKBUF_X2 inst_19073 ( .A(net_18920), .Z(net_18921) );
CLKBUF_X2 inst_14827 ( .A(net_14674), .Z(net_14675) );
CLKBUF_X2 inst_11324 ( .A(net_9364), .Z(net_11172) );
CLKBUF_X2 inst_15799 ( .A(net_12898), .Z(net_15647) );
CLKBUF_X2 inst_10696 ( .A(net_9710), .Z(net_10544) );
CLKBUF_X2 inst_13150 ( .A(net_12997), .Z(net_12998) );
SDFF_X2 inst_596 ( .SI(net_8389), .Q(net_8389), .SE(net_3969), .D(net_3958), .CK(net_10008) );
SDFFR_X1 inst_2771 ( .D(net_7378), .Q(net_7275), .SI(net_1956), .SE(net_1327), .CK(net_14663), .RN(x6501) );
AOI221_X2 inst_8835 ( .B1(net_8068), .C1(net_7864), .B2(net_6107), .ZN(net_6019), .C2(net_4400), .A(net_4294) );
NAND2_X2 inst_4687 ( .ZN(net_2011), .A1(net_2010), .A2(net_2007) );
CLKBUF_X2 inst_9245 ( .A(net_9092), .Z(net_9093) );
SDFF_X2 inst_1705 ( .SI(net_7847), .Q(net_7847), .D(net_2658), .SE(net_2558), .CK(net_15258) );
CLKBUF_X2 inst_11286 ( .A(net_10803), .Z(net_11134) );
NAND2_X2 inst_4664 ( .ZN(net_2447), .A2(net_2022), .A1(net_1744) );
CLKBUF_X2 inst_17388 ( .A(net_13756), .Z(net_17236) );
CLKBUF_X2 inst_14601 ( .A(net_14448), .Z(net_14449) );
MUX2_X2 inst_5003 ( .A(net_9036), .B(net_3990), .Z(net_3956), .S(net_622) );
CLKBUF_X2 inst_15841 ( .A(net_15688), .Z(net_15689) );
CLKBUF_X2 inst_12215 ( .A(net_10316), .Z(net_12063) );
CLKBUF_X2 inst_15454 ( .A(net_15301), .Z(net_15302) );
INV_X4 inst_5798 ( .A(net_6395), .ZN(net_2232) );
NOR3_X2 inst_3253 ( .A3(net_6179), .ZN(net_5689), .A1(net_5688), .A2(net_1366) );
INV_X4 inst_5321 ( .A(net_3162), .ZN(net_2528) );
CLKBUF_X2 inst_16378 ( .A(net_13477), .Z(net_16226) );
CLKBUF_X2 inst_14250 ( .A(net_14097), .Z(net_14098) );
NAND2_X2 inst_4596 ( .ZN(net_2778), .A1(net_2777), .A2(net_2775) );
AOI211_X2 inst_9013 ( .A(net_4924), .ZN(net_4838), .C1(net_4837), .C2(net_4836), .B(net_4821) );
AOI22_X2 inst_8427 ( .B1(net_6597), .A1(net_6564), .A2(net_6257), .B2(net_6110), .ZN(net_3514) );
CLKBUF_X2 inst_18316 ( .A(net_9372), .Z(net_18164) );
SDFF_X2 inst_637 ( .SI(net_8551), .Q(net_8551), .SE(net_3979), .D(net_3950), .CK(net_11001) );
CLKBUF_X2 inst_18649 ( .A(net_18496), .Z(net_18497) );
CLKBUF_X2 inst_13572 ( .A(net_13419), .Z(net_13420) );
CLKBUF_X2 inst_17211 ( .A(net_17058), .Z(net_17059) );
CLKBUF_X2 inst_18834 ( .A(net_18681), .Z(net_18682) );
CLKBUF_X2 inst_16024 ( .A(net_13497), .Z(net_15872) );
CLKBUF_X2 inst_13148 ( .A(net_12995), .Z(net_12996) );
DFFR_X2 inst_7033 ( .QN(net_7491), .D(net_5041), .CK(net_17258), .RN(x6501) );
CLKBUF_X2 inst_18496 ( .A(net_18343), .Z(net_18344) );
CLKBUF_X2 inst_15787 ( .A(net_13204), .Z(net_15635) );
AOI22_X2 inst_8152 ( .B2(net_8018), .A1(net_7984), .B1(net_6102), .A2(net_6097), .ZN(net_4000) );
CLKBUF_X2 inst_10159 ( .A(net_9784), .Z(net_10007) );
NAND2_X2 inst_4762 ( .ZN(net_1714), .A2(net_1379), .A1(net_897) );
XNOR2_X2 inst_164 ( .ZN(net_1839), .A(net_1572), .B(net_1552) );
AOI22_X2 inst_8534 ( .B1(net_6658), .A1(net_6625), .A2(net_6213), .B2(net_6138), .ZN(net_3406) );
AOI22_X2 inst_8467 ( .B1(net_6606), .A1(net_6573), .A2(net_6257), .B2(net_6110), .ZN(net_3473) );
SDFFR_X2 inst_2305 ( .SI(net_7408), .SE(net_2260), .Q(net_345), .D(net_345), .CK(net_9374), .RN(x6501) );
CLKBUF_X2 inst_10079 ( .A(net_9926), .Z(net_9927) );
SDFFR_X2 inst_2150 ( .Q(net_8273), .D(net_8273), .SI(net_3241), .SE(net_2996), .CK(net_18452), .RN(x6501) );
CLKBUF_X2 inst_10930 ( .A(net_10777), .Z(net_10778) );
CLKBUF_X2 inst_9770 ( .A(net_9617), .Z(net_9618) );
SDFF_X2 inst_946 ( .SI(net_7329), .Q(net_6703), .D(net_6703), .SE(net_3125), .CK(net_11654) );
SDFFR_X2 inst_2260 ( .SE(net_2801), .D(net_2760), .SI(net_206), .Q(net_206), .CK(net_14982), .RN(x6501) );
CLKBUF_X2 inst_18804 ( .A(net_12580), .Z(net_18652) );
AOI22_X2 inst_8141 ( .B1(net_8085), .A1(net_7745), .B2(net_6108), .A2(net_6096), .ZN(net_4010) );
CLKBUF_X2 inst_13276 ( .A(net_13123), .Z(net_13124) );
CLKBUF_X2 inst_19048 ( .A(net_10269), .Z(net_18896) );
CLKBUF_X2 inst_11700 ( .A(net_11547), .Z(net_11548) );
NAND2_X2 inst_4625 ( .ZN(net_2581), .A2(net_2471), .A1(net_2160) );
DFFS_X1 inst_6951 ( .D(net_6145), .CK(net_13616), .SN(x6501), .Q(x785) );
NAND3_X2 inst_3922 ( .ZN(net_5616), .A1(net_5545), .A3(net_5479), .A2(net_5303) );
SDFF_X2 inst_2053 ( .SI(net_7800), .Q(net_7800), .D(net_2715), .SE(net_2459), .CK(net_16790) );
CLKBUF_X2 inst_10539 ( .A(net_10386), .Z(net_10387) );
CLKBUF_X2 inst_10038 ( .A(net_9178), .Z(net_9886) );
SDFF_X2 inst_1325 ( .SI(net_7697), .Q(net_7697), .SE(net_2714), .D(net_2639), .CK(net_16512) );
CLKBUF_X2 inst_19018 ( .A(net_15232), .Z(net_18866) );
AOI221_X2 inst_8859 ( .ZN(net_2988), .B2(net_2967), .C2(net_2943), .A(net_2839), .C1(net_1715), .B1(net_870) );
CLKBUF_X2 inst_17861 ( .A(net_13543), .Z(net_17709) );
CLKBUF_X2 inst_13503 ( .A(net_13350), .Z(net_13351) );
CLKBUF_X2 inst_16684 ( .A(net_16531), .Z(net_16532) );
DFFS_X2 inst_6873 ( .QN(net_8294), .D(net_3968), .CK(net_11199), .SN(x6501) );
CLKBUF_X2 inst_14087 ( .A(net_13934), .Z(net_13935) );
NOR3_X2 inst_3312 ( .A2(net_9049), .ZN(net_3949), .A1(net_1458), .A3(net_622) );
CLKBUF_X2 inst_15432 ( .A(net_15279), .Z(net_15280) );
AND2_X2 inst_9207 ( .ZN(net_1339), .A1(net_1186), .A2(net_846) );
CLKBUF_X2 inst_17138 ( .A(net_16985), .Z(net_16986) );
CLKBUF_X2 inst_12143 ( .A(net_9465), .Z(net_11991) );
SDFF_X2 inst_1235 ( .Q(net_7810), .D(net_7810), .SE(net_2730), .SI(net_2709), .CK(net_15857) );
CLKBUF_X2 inst_16948 ( .A(net_14697), .Z(net_16796) );
CLKBUF_X2 inst_16760 ( .A(net_14664), .Z(net_16608) );
CLKBUF_X2 inst_15015 ( .A(net_12646), .Z(net_14863) );
CLKBUF_X2 inst_14107 ( .A(net_13954), .Z(net_13955) );
CLKBUF_X2 inst_13143 ( .A(net_12990), .Z(net_12991) );
CLKBUF_X2 inst_16115 ( .A(net_11563), .Z(net_15963) );
NAND4_X2 inst_3626 ( .A4(net_6792), .ZN(net_5814), .A2(net_2028), .A3(net_1062), .A1(net_1058) );
NAND2_X4 inst_4036 ( .ZN(net_4928), .A2(net_4800), .A1(net_2580) );
INV_X4 inst_5244 ( .A(net_2028), .ZN(net_1912) );
CLKBUF_X2 inst_19068 ( .A(net_18915), .Z(net_18916) );
CLKBUF_X2 inst_14942 ( .A(net_14789), .Z(net_14790) );
CLKBUF_X2 inst_13457 ( .A(net_13304), .Z(net_13305) );
CLKBUF_X2 inst_18572 ( .A(net_18419), .Z(net_18420) );
SDFF_X2 inst_1600 ( .Q(net_8135), .D(net_8135), .SI(net_2749), .SE(net_2541), .CK(net_17135) );
OR2_X4 inst_2850 ( .A1(net_9054), .A2(net_3161), .ZN(net_2532) );
CLKBUF_X2 inst_14884 ( .A(net_14731), .Z(net_14732) );
CLKBUF_X2 inst_14268 ( .A(net_14115), .Z(net_14116) );
INV_X4 inst_5163 ( .ZN(net_3177), .A(net_3157) );
CLKBUF_X2 inst_9590 ( .A(net_9380), .Z(net_9438) );
SDFF_X2 inst_849 ( .SI(net_8661), .Q(net_8661), .D(net_3951), .SE(net_3885), .CK(net_12860) );
DFFR_X1 inst_7393 ( .QN(net_6300), .D(net_5854), .CK(net_16775), .RN(x6501) );
CLKBUF_X2 inst_16998 ( .A(net_14287), .Z(net_16846) );
XOR2_X2 inst_3 ( .Z(net_3207), .A(net_2996), .B(net_2989) );
CLKBUF_X2 inst_14517 ( .A(net_14364), .Z(net_14365) );
OAI21_X2 inst_3060 ( .B2(net_8244), .B1(net_4850), .ZN(net_4747), .A(net_2603) );
INV_X4 inst_5812 ( .A(net_7396), .ZN(net_1779) );
CLKBUF_X2 inst_10041 ( .A(net_9888), .Z(net_9889) );
SDFF_X2 inst_566 ( .Q(net_8829), .D(net_8829), .SE(net_3964), .SI(net_3959), .CK(net_13200) );
SDFF_X2 inst_1399 ( .Q(net_8204), .D(net_8204), .SI(net_2717), .SE(net_2561), .CK(net_14183) );
CLKBUF_X2 inst_19180 ( .A(net_19027), .Z(net_19028) );
CLKBUF_X2 inst_12301 ( .A(net_12148), .Z(net_12149) );
CLKBUF_X2 inst_10613 ( .A(net_9614), .Z(net_10461) );
NAND2_X2 inst_4357 ( .A1(net_7082), .A2(net_5164), .ZN(net_5100) );
CLKBUF_X2 inst_16456 ( .A(net_16303), .Z(net_16304) );
NAND2_X2 inst_4327 ( .A1(net_7100), .A2(net_5164), .ZN(net_5130) );
CLKBUF_X2 inst_16189 ( .A(net_16036), .Z(net_16037) );
CLKBUF_X2 inst_11375 ( .A(net_10773), .Z(net_11223) );
CLKBUF_X2 inst_10419 ( .A(net_10266), .Z(net_10267) );
SDFFR_X2 inst_2333 ( .SI(net_7373), .SE(net_2732), .D(net_1052), .QN(net_148), .CK(net_16129), .RN(x6501) );
CLKBUF_X2 inst_14844 ( .A(net_14691), .Z(net_14692) );
CLKBUF_X2 inst_15291 ( .A(net_15138), .Z(net_15139) );
DFFR_X2 inst_7047 ( .QN(net_7498), .D(net_4842), .CK(net_14491), .RN(x6501) );
CLKBUF_X2 inst_11345 ( .A(net_11192), .Z(net_11193) );
INV_X4 inst_5928 ( .A(net_6816), .ZN(net_4621) );
INV_X8 inst_5056 ( .A(net_6261), .ZN(net_6260) );
INV_X4 inst_5370 ( .ZN(net_1132), .A(net_1131) );
SDFF_X2 inst_1732 ( .Q(net_7987), .D(net_7987), .SI(net_2706), .SE(net_2542), .CK(net_15238) );
DFFR_X2 inst_7256 ( .Q(net_7485), .D(net_296), .CK(net_13458), .RN(x6501) );
CLKBUF_X2 inst_18697 ( .A(net_18544), .Z(net_18545) );
INV_X4 inst_6119 ( .A(net_7235), .ZN(net_1807) );
CLKBUF_X2 inst_15461 ( .A(net_15308), .Z(net_15309) );
INV_X2 inst_6269 ( .A(net_8230), .ZN(net_4627) );
CLKBUF_X2 inst_13247 ( .A(net_12033), .Z(net_13095) );
CLKBUF_X2 inst_9481 ( .A(net_9328), .Z(net_9329) );
INV_X4 inst_5858 ( .A(net_8257), .ZN(net_1211) );
OAI21_X2 inst_3069 ( .B2(net_6444), .B1(net_4362), .ZN(net_4312), .A(net_2956) );
NAND4_X2 inst_3631 ( .ZN(net_5537), .A4(net_5275), .A3(net_4702), .A1(net_4542), .A2(net_4541) );
SDFF_X2 inst_1101 ( .D(net_7312), .SI(net_6521), .Q(net_6521), .SE(net_3086), .CK(net_12006) );
AOI222_X1 inst_8596 ( .B2(net_6773), .B1(net_5835), .C2(net_5832), .ZN(net_5831), .A2(net_5830), .A1(net_3268), .C1(x2908) );
CLKBUF_X2 inst_17712 ( .A(net_17101), .Z(net_17560) );
INV_X1 inst_6652 ( .ZN(net_2171), .A(net_2170) );
OAI221_X2 inst_2950 ( .B1(net_7571), .B2(net_4971), .ZN(net_4959), .C1(net_4928), .C2(net_4628), .A(net_2917) );
AOI22_X2 inst_8584 ( .B2(net_6320), .ZN(net_1788), .A2(net_1253), .B1(net_1252), .A1(x4347) );
CLKBUF_X2 inst_15777 ( .A(net_15595), .Z(net_15625) );
CLKBUF_X2 inst_17673 ( .A(net_17520), .Z(net_17521) );
CLKBUF_X2 inst_12013 ( .A(net_11860), .Z(net_11861) );
CLKBUF_X2 inst_15572 ( .A(net_15419), .Z(net_15420) );
SDFFR_X2 inst_2451 ( .D(net_3236), .SE(net_2678), .SI(net_420), .Q(net_420), .CK(net_17271), .RN(x6501) );
CLKBUF_X2 inst_16326 ( .A(net_16173), .Z(net_16174) );
SDFF_X2 inst_1202 ( .D(net_7300), .SI(net_6997), .Q(net_6997), .SE(net_6283), .CK(net_15918) );
CLKBUF_X2 inst_15106 ( .A(net_14953), .Z(net_14954) );
DFFR_X2 inst_7020 ( .QN(net_6306), .D(net_5711), .CK(net_14217), .RN(x6501) );
SDFFR_X2 inst_2227 ( .Q(net_7474), .D(net_7474), .SE(net_2863), .CK(net_12178), .SI(x13396), .RN(x6501) );
SDFF_X2 inst_660 ( .Q(net_8434), .D(net_8434), .SI(net_3975), .SE(net_3934), .CK(net_10253) );
SDFFR_X2 inst_2490 ( .Q(net_8983), .D(net_8983), .SI(net_2616), .SE(net_2562), .CK(net_17269), .RN(x6501) );
CLKBUF_X2 inst_14526 ( .A(net_14373), .Z(net_14374) );
CLKBUF_X2 inst_10150 ( .A(net_9997), .Z(net_9998) );
SDFF_X2 inst_1576 ( .Q(net_8026), .D(net_8026), .SI(net_2575), .SE(net_2545), .CK(net_16044) );
CLKBUF_X2 inst_16712 ( .A(net_16559), .Z(net_16560) );
CLKBUF_X2 inst_11532 ( .A(net_10636), .Z(net_11380) );
INV_X4 inst_5642 ( .A(net_6422), .ZN(net_1830) );
CLKBUF_X2 inst_16397 ( .A(net_16244), .Z(net_16245) );
DFFR_X1 inst_7459 ( .QN(net_6795), .D(net_6192), .CK(net_9595), .RN(x6501) );
CLKBUF_X2 inst_11898 ( .A(net_11745), .Z(net_11746) );
AOI22_X2 inst_8390 ( .B1(net_8858), .A1(net_8303), .B2(net_6252), .A2(net_4345), .ZN(net_3659) );
CLKBUF_X2 inst_17141 ( .A(net_16988), .Z(net_16989) );
INV_X1 inst_6659 ( .A(net_6198), .ZN(net_6196) );
CLKBUF_X2 inst_18859 ( .A(net_18706), .Z(net_18707) );
AOI22_X2 inst_7828 ( .A2(net_5535), .B2(net_5260), .ZN(net_4693), .B1(net_2968), .A1(net_453) );
NAND2_X2 inst_4368 ( .A1(net_7153), .A2(net_5166), .ZN(net_5089) );
CLKBUF_X2 inst_10331 ( .A(net_10178), .Z(net_10179) );
CLKBUF_X2 inst_11137 ( .A(net_10984), .Z(net_10985) );
CLKBUF_X2 inst_17604 ( .A(net_17451), .Z(net_17452) );
SDFF_X2 inst_1147 ( .SI(net_7328), .Q(net_6603), .D(net_6603), .SE(net_3069), .CK(net_11750) );
SDFF_X2 inst_1768 ( .D(net_7297), .SI(net_6874), .Q(net_6874), .SE(net_6282), .CK(net_15427) );
CLKBUF_X2 inst_18308 ( .A(net_18155), .Z(net_18156) );
INV_X2 inst_6410 ( .A(net_1333), .ZN(net_1064) );
CLKBUF_X2 inst_12865 ( .A(net_12712), .Z(net_12713) );
OAI22_X2 inst_2917 ( .ZN(net_3539), .A2(net_3538), .B2(net_3537), .A1(net_3162), .B1(net_746) );
CLKBUF_X2 inst_18953 ( .A(net_18800), .Z(net_18801) );
SDFF_X2 inst_1408 ( .SI(net_7283), .Q(net_7140), .D(net_7140), .SE(net_6279), .CK(net_16240) );
CLKBUF_X2 inst_13563 ( .A(net_13410), .Z(net_13411) );
SDFF_X2 inst_1889 ( .D(net_7270), .SI(net_6967), .Q(net_6967), .SE(net_6283), .CK(net_14333) );
SDFF_X2 inst_2011 ( .SI(net_7804), .Q(net_7804), .D(net_2656), .SE(net_2459), .CK(net_14384) );
CLKBUF_X2 inst_13495 ( .A(net_11750), .Z(net_13343) );
SDFF_X2 inst_1761 ( .SI(net_7759), .Q(net_7759), .D(net_2713), .SE(net_2560), .CK(net_16468) );
CLKBUF_X2 inst_16000 ( .A(net_15847), .Z(net_15848) );
INV_X2 inst_6582 ( .A(net_7428), .ZN(net_480) );
CLKBUF_X2 inst_9418 ( .A(net_9265), .Z(net_9266) );
INV_X4 inst_5474 ( .A(net_2876), .ZN(net_745) );
XOR2_X1 inst_84 ( .Z(net_2985), .A(net_2821), .B(x3028) );
INV_X4 inst_5974 ( .A(net_8898), .ZN(net_1074) );
XNOR2_X2 inst_173 ( .B(net_2389), .ZN(net_1791), .A(net_1790) );
INV_X4 inst_5568 ( .A(net_7372), .ZN(net_1226) );
INV_X4 inst_5821 ( .A(net_7352), .ZN(net_737) );
DFFR_X2 inst_7187 ( .QN(net_7362), .D(net_2495), .CK(net_11833), .RN(x6501) );
INV_X4 inst_5713 ( .ZN(net_916), .A(net_395) );
CLKBUF_X2 inst_10493 ( .A(net_10340), .Z(net_10341) );
AOI221_X4 inst_8723 ( .B1(net_8816), .C1(net_8335), .C2(net_6265), .B2(net_6253), .ZN(net_4343), .A(net_4256) );
CLKBUF_X2 inst_13047 ( .A(net_12894), .Z(net_12895) );
SDFF_X2 inst_1943 ( .SI(net_8077), .Q(net_8077), .D(net_2703), .SE(net_2508), .CK(net_13994) );
AOI22_X2 inst_7847 ( .B2(net_5609), .A2(net_5595), .ZN(net_4661), .B1(net_351), .A1(net_307) );
INV_X4 inst_5573 ( .A(net_5980), .ZN(x3762) );
CLKBUF_X2 inst_18598 ( .A(net_18445), .Z(net_18446) );
SDFF_X2 inst_1531 ( .Q(net_7877), .D(net_7877), .SI(net_2655), .SE(net_2543), .CK(net_15445) );
DFFR_X2 inst_7083 ( .QN(net_7664), .D(net_3893), .CK(net_12678), .RN(x6501) );
CLKBUF_X2 inst_11706 ( .A(net_10446), .Z(net_11554) );
CLKBUF_X2 inst_15075 ( .A(net_14922), .Z(net_14923) );
OAI22_X2 inst_2922 ( .A2(net_3064), .ZN(net_2987), .B2(net_2834), .B1(net_2206), .A1(net_1165) );
CLKBUF_X2 inst_11831 ( .A(net_9293), .Z(net_11679) );
CLKBUF_X2 inst_11649 ( .A(net_11496), .Z(net_11497) );
CLKBUF_X2 inst_10410 ( .A(net_10257), .Z(net_10258) );
CLKBUF_X2 inst_18551 ( .A(net_15702), .Z(net_18399) );
CLKBUF_X2 inst_18682 ( .A(net_11878), .Z(net_18530) );
CLKBUF_X2 inst_16036 ( .A(net_15883), .Z(net_15884) );
SDFF_X2 inst_1037 ( .SI(net_7323), .Q(net_6730), .D(net_6730), .SE(net_3124), .CK(net_9137) );
AOI22_X2 inst_7777 ( .B1(net_6967), .A1(net_6927), .A2(net_5443), .B2(net_5442), .ZN(net_5295) );
AOI222_X1 inst_8652 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3914), .B1(net_3100), .C1(net_3098), .A1(x13761) );
NOR2_X2 inst_3596 ( .ZN(net_3328), .A1(net_1150), .A2(net_1074) );
SDFF_X2 inst_1250 ( .SI(net_7695), .Q(net_7695), .SE(net_2714), .D(net_2711), .CK(net_14188) );
DFFR_X2 inst_7071 ( .QN(net_7415), .D(net_4204), .CK(net_12298), .RN(x6501) );
CLKBUF_X2 inst_10240 ( .A(net_9997), .Z(net_10088) );
CLKBUF_X2 inst_19028 ( .A(net_18875), .Z(net_18876) );
SDFF_X2 inst_1979 ( .D(net_7294), .SI(net_6911), .Q(net_6911), .SE(net_6284), .CK(net_17655) );
SDFF_X2 inst_364 ( .SI(net_8301), .Q(net_8301), .SE(net_3978), .D(net_3938), .CK(net_12480) );
CLKBUF_X2 inst_11586 ( .A(net_11433), .Z(net_11434) );
CLKBUF_X2 inst_9253 ( .A(net_9093), .Z(net_9101) );
CLKBUF_X2 inst_9283 ( .A(net_9130), .Z(net_9131) );
OAI21_X2 inst_2997 ( .B2(net_5902), .ZN(net_5896), .A(net_5827), .B1(net_781) );
NAND2_X2 inst_4712 ( .ZN(net_2585), .A1(net_1877), .A2(net_1586) );
SDFF_X2 inst_411 ( .SI(net_8325), .Q(net_8325), .SE(net_3978), .D(net_3953), .CK(net_10298) );
AND2_X4 inst_9055 ( .ZN(net_6266), .A1(net_3352), .A2(net_3351) );
CLKBUF_X2 inst_10380 ( .A(net_9565), .Z(net_10228) );
NAND2_X4 inst_4026 ( .ZN(net_6143), .A2(net_6088), .A1(net_6087) );
CLKBUF_X2 inst_14722 ( .A(net_14569), .Z(net_14570) );
CLKBUF_X2 inst_14649 ( .A(net_9394), .Z(net_14497) );
CLKBUF_X2 inst_9395 ( .A(net_9137), .Z(net_9243) );
CLKBUF_X2 inst_11333 ( .A(net_10649), .Z(net_11181) );
CLKBUF_X2 inst_10668 ( .A(net_10515), .Z(net_10516) );
CLKBUF_X2 inst_11010 ( .A(net_10857), .Z(net_10858) );
NAND2_X2 inst_4382 ( .A1(net_7077), .A2(net_5162), .ZN(net_5075) );
CLKBUF_X2 inst_10908 ( .A(net_10755), .Z(net_10756) );
CLKBUF_X2 inst_14426 ( .A(net_14273), .Z(net_14274) );
CLKBUF_X2 inst_17391 ( .A(net_17238), .Z(net_17239) );
CLKBUF_X2 inst_13480 ( .A(net_13327), .Z(net_13328) );
CLKBUF_X2 inst_17941 ( .A(net_15972), .Z(net_17789) );
AOI221_X4 inst_8708 ( .C1(net_8200), .B1(net_7690), .C2(net_6099), .ZN(net_6039), .B2(net_4399), .A(net_4298) );
CLKBUF_X2 inst_15400 ( .A(net_13874), .Z(net_15248) );
CLKBUF_X2 inst_13297 ( .A(net_11821), .Z(net_13145) );
CLKBUF_X2 inst_14020 ( .A(net_12089), .Z(net_13868) );
CLKBUF_X2 inst_9874 ( .A(net_9721), .Z(net_9722) );
INV_X4 inst_5538 ( .ZN(net_875), .A(net_652) );
XOR2_X2 inst_61 ( .B(net_1877), .A(net_1778), .Z(net_942) );
XNOR2_X2 inst_203 ( .ZN(net_1540), .A(net_926), .B(net_924) );
INV_X4 inst_5834 ( .A(net_8896), .ZN(net_913) );
CLKBUF_X2 inst_14077 ( .A(net_13924), .Z(net_13925) );
SDFF_X2 inst_1139 ( .D(net_7318), .SI(net_6560), .Q(net_6560), .SE(net_3070), .CK(net_9909) );
CLKBUF_X2 inst_10597 ( .A(net_9846), .Z(net_10445) );
AOI221_X2 inst_8852 ( .B1(net_8580), .C1(net_8469), .C2(net_6263), .B2(net_6262), .ZN(net_6225), .A(net_4251) );
NAND2_X2 inst_4507 ( .A2(net_6272), .ZN(net_4356), .A1(net_4355) );
CLKBUF_X2 inst_17381 ( .A(net_12826), .Z(net_17229) );
CLKBUF_X2 inst_14558 ( .A(net_14405), .Z(net_14406) );
CLKBUF_X2 inst_9968 ( .A(net_9815), .Z(net_9816) );
CLKBUF_X2 inst_14669 ( .A(net_14516), .Z(net_14517) );
INV_X2 inst_6607 ( .A(net_6169), .ZN(net_6166) );
SDFF_X2 inst_456 ( .SI(net_8458), .Q(net_8458), .SE(net_3983), .D(net_3966), .CK(net_13280) );
SDFF_X2 inst_832 ( .SI(net_8641), .Q(net_8641), .D(net_3962), .SE(net_3885), .CK(net_10144) );
AOI22_X2 inst_8102 ( .B1(net_8076), .A1(net_7872), .B2(net_6107), .A2(net_4400), .ZN(net_4046) );
XNOR2_X2 inst_275 ( .ZN(net_1034), .A(net_1033), .B(net_198) );
CLKBUF_X2 inst_11492 ( .A(net_11339), .Z(net_11340) );
NAND4_X2 inst_3728 ( .ZN(net_4302), .A1(net_4148), .A2(net_4147), .A3(net_4146), .A4(net_4145) );
CLKBUF_X2 inst_11576 ( .A(net_11423), .Z(net_11424) );
SDFFR_X2 inst_2416 ( .D(net_2688), .SE(net_2313), .SI(net_460), .Q(net_460), .CK(net_16916), .RN(x6501) );
CLKBUF_X2 inst_17239 ( .A(net_17086), .Z(net_17087) );
NAND4_X2 inst_3812 ( .ZN(net_3614), .A1(net_3439), .A2(net_3438), .A3(net_3437), .A4(net_3436) );
CLKBUF_X2 inst_17069 ( .A(net_14569), .Z(net_16917) );
AOI22_X2 inst_7879 ( .A2(net_5538), .ZN(net_4556), .B2(net_4555), .B1(net_1805), .A1(net_432) );
NAND3_X2 inst_3959 ( .ZN(net_3072), .A2(net_2946), .A3(net_2945), .A1(net_2899) );
CLKBUF_X2 inst_9839 ( .A(net_9686), .Z(net_9687) );
NAND2_X2 inst_4518 ( .ZN(net_4837), .A2(net_4554), .A1(net_1600) );
CLKBUF_X2 inst_11185 ( .A(net_10014), .Z(net_11033) );
CLKBUF_X2 inst_15415 ( .A(net_9074), .Z(net_15263) );
CLKBUF_X2 inst_10348 ( .A(net_10195), .Z(net_10196) );
CLKBUF_X2 inst_9726 ( .A(net_9573), .Z(net_9574) );
DFF_X1 inst_6832 ( .Q(net_6452), .D(net_3616), .CK(net_15164) );
CLKBUF_X2 inst_14234 ( .A(net_9642), .Z(net_14082) );
AOI22_X2 inst_7958 ( .A1(net_7955), .B1(net_7785), .A2(net_6092), .B2(net_6091), .ZN(net_4169) );
CLKBUF_X2 inst_11237 ( .A(net_11084), .Z(net_11085) );
OAI21_X2 inst_3166 ( .ZN(net_1609), .A(net_1608), .B2(net_1607), .B1(net_542) );
CLKBUF_X2 inst_18131 ( .A(net_14806), .Z(net_17979) );
CLKBUF_X2 inst_14218 ( .A(net_14065), .Z(net_14066) );
DFFR_X1 inst_7452 ( .QN(net_8935), .D(net_4747), .CK(net_14581), .RN(x6501) );
CLKBUF_X2 inst_13807 ( .A(net_12919), .Z(net_13655) );
NAND4_X2 inst_3656 ( .A4(net_6006), .A1(net_6005), .ZN(net_4609), .A2(net_4156), .A3(net_4155) );
CLKBUF_X2 inst_12497 ( .A(net_12344), .Z(net_12345) );
SDFFR_X2 inst_2237 ( .Q(net_7461), .D(net_7461), .SE(net_2863), .CK(net_10625), .SI(x13501), .RN(x6501) );
AND2_X2 inst_9155 ( .ZN(net_2875), .A2(net_2874), .A1(net_1071) );
CLKBUF_X2 inst_14905 ( .A(net_14752), .Z(net_14753) );
CLKBUF_X2 inst_14570 ( .A(net_14417), .Z(net_14418) );
DFF_X1 inst_6834 ( .Q(net_6454), .D(net_3614), .CK(net_15156) );
CLKBUF_X2 inst_18175 ( .A(net_16340), .Z(net_18023) );
CLKBUF_X2 inst_18407 ( .A(net_15821), .Z(net_18255) );
CLKBUF_X2 inst_10701 ( .A(net_9474), .Z(net_10549) );
OR2_X4 inst_2827 ( .ZN(net_3571), .A1(net_3570), .A2(net_3527) );
AND2_X4 inst_9062 ( .A1(net_3318), .A2(net_3305), .ZN(net_3302) );
SDFFR_X2 inst_2448 ( .D(net_3051), .SE(net_2683), .SI(net_415), .Q(net_415), .CK(net_17275), .RN(x6501) );
CLKBUF_X2 inst_17146 ( .A(net_16993), .Z(net_16994) );
SDFFR_X2 inst_2541 ( .QN(net_6364), .SE(net_2147), .D(net_2143), .SI(net_1950), .CK(net_14755), .RN(x6501) );
CLKBUF_X2 inst_17525 ( .A(net_10674), .Z(net_17373) );
SDFF_X2 inst_1693 ( .Q(net_8147), .D(net_8147), .SI(net_2585), .SE(net_2538), .CK(net_18524) );
NOR3_X2 inst_3306 ( .A1(net_2731), .A2(net_2698), .ZN(net_1660), .A3(net_1257) );
SDFF_X2 inst_1020 ( .SI(net_7335), .Q(net_6676), .D(net_6676), .SE(net_3126), .CK(net_9763) );
CLKBUF_X2 inst_11007 ( .A(net_9326), .Z(net_10855) );
CLKBUF_X2 inst_17959 ( .A(net_17806), .Z(net_17807) );
CLKBUF_X2 inst_11057 ( .A(net_10904), .Z(net_10905) );
CLKBUF_X2 inst_13886 ( .A(net_13733), .Z(net_13734) );
CLKBUF_X2 inst_16298 ( .A(net_16145), .Z(net_16146) );
NAND3_X2 inst_3952 ( .ZN(net_3336), .A3(net_3308), .A1(net_3242), .A2(net_1151) );
CLKBUF_X2 inst_12084 ( .A(net_11931), .Z(net_11932) );
NOR2_X2 inst_3588 ( .A2(net_8895), .ZN(net_3245), .A1(net_913) );
CLKBUF_X2 inst_15120 ( .A(net_12199), .Z(net_14968) );
INV_X4 inst_5559 ( .ZN(net_1480), .A(net_625) );
SDFF_X2 inst_1096 ( .D(net_7322), .SI(net_6531), .Q(net_6531), .SE(net_3086), .CK(net_9151) );
CLKBUF_X2 inst_16336 ( .A(net_11102), .Z(net_16184) );
NAND2_X2 inst_4552 ( .A1(net_6255), .ZN(net_3526), .A2(net_3304) );
CLKBUF_X2 inst_9260 ( .A(net_9099), .Z(net_9108) );
INV_X4 inst_5637 ( .A(net_7479), .ZN(net_3127) );
SDFF_X2 inst_1839 ( .D(net_7280), .SI(net_6897), .Q(net_6897), .SE(net_6284), .CK(net_18999) );
CLKBUF_X2 inst_14708 ( .A(net_12741), .Z(net_14556) );
CLKBUF_X2 inst_18332 ( .A(net_13978), .Z(net_18180) );
AOI22_X2 inst_8041 ( .B1(net_8034), .A1(net_8000), .B2(net_6102), .A2(net_6097), .ZN(net_4098) );
CLKBUF_X2 inst_13095 ( .A(net_12942), .Z(net_12943) );
SDFF_X2 inst_725 ( .SI(net_8509), .Q(net_8509), .D(net_3941), .SE(net_3884), .CK(net_10343) );
CLKBUF_X2 inst_12840 ( .A(net_12687), .Z(net_12688) );
INV_X2 inst_6326 ( .ZN(net_3264), .A(net_3263) );
SDFF_X2 inst_1337 ( .Q(net_7947), .D(net_7947), .SE(net_2755), .SI(net_2659), .CK(net_18076) );
CLKBUF_X2 inst_18181 ( .A(net_18028), .Z(net_18029) );
INV_X4 inst_5375 ( .ZN(net_1124), .A(x3485) );
OAI21_X2 inst_3096 ( .B1(net_6117), .ZN(net_2780), .B2(net_2487), .A(net_2211) );
CLKBUF_X2 inst_15532 ( .A(net_15379), .Z(net_15380) );
OAI21_X2 inst_3015 ( .A(net_6249), .B1(net_6179), .ZN(net_5273), .B2(net_5272) );
CLKBUF_X2 inst_11618 ( .A(net_11465), .Z(net_11466) );
SDFFR_X2 inst_2441 ( .D(net_3239), .SE(net_2757), .SI(net_425), .Q(net_425), .CK(net_17276), .RN(x6501) );
CLKBUF_X2 inst_17288 ( .A(net_9758), .Z(net_17136) );
CLKBUF_X2 inst_16264 ( .A(net_16111), .Z(net_16112) );
CLKBUF_X2 inst_11945 ( .A(net_11792), .Z(net_11793) );
CLKBUF_X2 inst_9714 ( .A(net_9561), .Z(net_9562) );
DFFR_X1 inst_7427 ( .QN(net_8910), .D(net_4860), .CK(net_14854), .RN(x6501) );
SDFF_X2 inst_878 ( .Q(net_8590), .D(net_8590), .SI(net_3939), .SE(net_3878), .CK(net_12493) );
CLKBUF_X2 inst_17099 ( .A(net_13894), .Z(net_16947) );
MUX2_X2 inst_4959 ( .A(net_7377), .S(net_2376), .Z(net_2364), .B(net_828) );
CLKBUF_X2 inst_18707 ( .A(net_18554), .Z(net_18555) );
CLKBUF_X2 inst_13442 ( .A(net_13289), .Z(net_13290) );
DFF_X1 inst_6782 ( .Q(net_7531), .D(net_4588), .CK(net_11966) );
SDFF_X2 inst_1926 ( .SI(net_8053), .Q(net_8053), .D(net_2573), .SE(net_2508), .CK(net_18030) );
NAND2_X2 inst_4351 ( .A1(net_7108), .A2(net_5164), .ZN(net_5106) );
CLKBUF_X2 inst_17683 ( .A(net_17530), .Z(net_17531) );
CLKBUF_X2 inst_16908 ( .A(net_10579), .Z(net_16756) );
INV_X2 inst_6211 ( .ZN(net_5499), .A(net_5385) );
CLKBUF_X2 inst_12761 ( .A(net_12608), .Z(net_12609) );
INV_X2 inst_6383 ( .ZN(net_1332), .A(net_1331) );
SDFF_X2 inst_564 ( .Q(net_8827), .D(net_8827), .SE(net_3964), .SI(net_3945), .CK(net_13133) );
CLKBUF_X2 inst_12795 ( .A(net_12642), .Z(net_12643) );
CLKBUF_X2 inst_10262 ( .A(net_9842), .Z(net_10110) );
CLKBUF_X2 inst_16913 ( .A(net_16760), .Z(net_16761) );
CLKBUF_X2 inst_11210 ( .A(net_11057), .Z(net_11058) );
INV_X2 inst_6500 ( .A(net_7510), .ZN(net_541) );
SDFF_X2 inst_934 ( .SI(net_7341), .Q(net_6682), .D(net_6682), .SE(net_3126), .CK(net_11692) );
SDFF_X2 inst_1000 ( .D(net_7340), .SI(net_6648), .Q(net_6648), .SE(net_3123), .CK(net_11908) );
CLKBUF_X2 inst_17398 ( .A(net_17245), .Z(net_17246) );
CLKBUF_X2 inst_18606 ( .A(net_18453), .Z(net_18454) );
CLKBUF_X2 inst_18188 ( .A(net_18035), .Z(net_18036) );
SDFFR_X2 inst_2585 ( .D(net_7377), .QN(net_7237), .SI(net_1952), .SE(net_1379), .CK(net_14651), .RN(x6501) );
CLKBUF_X2 inst_12044 ( .A(net_10438), .Z(net_11892) );
SDFFR_X2 inst_2364 ( .SI(net_7378), .D(net_2724), .SE(net_2723), .QN(net_159), .CK(net_17815), .RN(x6501) );
NAND2_X2 inst_4299 ( .A1(net_7132), .A2(net_5166), .ZN(net_5158) );
CLKBUF_X2 inst_18502 ( .A(net_18349), .Z(net_18350) );
CLKBUF_X2 inst_11281 ( .A(net_9074), .Z(net_11129) );
SDFF_X2 inst_1882 ( .D(net_7292), .SI(net_6989), .Q(net_6989), .SE(net_6283), .CK(net_14875) );
CLKBUF_X2 inst_14510 ( .A(net_14357), .Z(net_14358) );
CLKBUF_X2 inst_13787 ( .A(net_10649), .Z(net_13635) );
CLKBUF_X2 inst_14482 ( .A(net_9812), .Z(net_14330) );
AOI22_X2 inst_7812 ( .A2(net_8239), .B2(net_6144), .A1(net_4764), .ZN(net_4752), .B1(net_4551) );
CLKBUF_X2 inst_17273 ( .A(net_17120), .Z(net_17121) );
AOI22_X2 inst_8441 ( .B1(net_6667), .A1(net_6634), .A2(net_6213), .B2(net_6138), .ZN(net_3500) );
AOI22_X2 inst_8218 ( .A1(net_8610), .B1(net_8425), .A2(net_3864), .B2(net_3863), .ZN(net_3818) );
INV_X2 inst_6578 ( .ZN(net_851), .A(net_228) );
CLKBUF_X2 inst_19174 ( .A(net_15651), .Z(net_19022) );
CLKBUF_X2 inst_16149 ( .A(net_14451), .Z(net_15997) );
CLKBUF_X2 inst_12849 ( .A(net_12696), .Z(net_12697) );
CLKBUF_X2 inst_17686 ( .A(net_17533), .Z(net_17534) );
INV_X4 inst_5531 ( .A(net_909), .ZN(net_659) );
INV_X4 inst_5397 ( .A(net_885), .ZN(x3485) );
SDFF_X2 inst_727 ( .SI(net_8483), .Q(net_8483), .D(net_3943), .SE(net_3884), .CK(net_13100) );
CLKBUF_X2 inst_11795 ( .A(net_11642), .Z(net_11643) );
NAND2_X2 inst_4804 ( .A2(net_7399), .ZN(net_1584), .A1(net_1087) );
CLKBUF_X2 inst_11686 ( .A(net_11533), .Z(net_11534) );
OR2_X2 inst_2874 ( .ZN(net_4413), .A1(net_4412), .A2(net_4411) );
INV_X2 inst_6485 ( .ZN(net_560), .A(net_386) );
NAND2_X2 inst_4607 ( .A2(net_6144), .ZN(net_2627), .A1(net_2626) );
SDFFR_X2 inst_2431 ( .SE(net_2748), .D(net_2672), .SI(net_435), .Q(net_435), .CK(net_14552), .RN(x6501) );
AOI221_X2 inst_8861 ( .ZN(net_3323), .B2(net_2244), .C1(net_2179), .C2(net_1998), .A(net_1892), .B1(net_1262) );
CLKBUF_X2 inst_12052 ( .A(net_11899), .Z(net_11900) );
CLKBUF_X2 inst_18713 ( .A(net_18560), .Z(net_18561) );
AOI22_X2 inst_8274 ( .B1(net_8765), .A1(net_8395), .A2(net_3867), .B2(net_3866), .ZN(net_3766) );
CLKBUF_X2 inst_16085 ( .A(net_15932), .Z(net_15933) );
SDFF_X2 inst_953 ( .SI(net_7340), .Q(net_6714), .D(net_6714), .SE(net_3125), .CK(net_11921) );
CLKBUF_X2 inst_16605 ( .A(net_16233), .Z(net_16453) );
CLKBUF_X2 inst_13674 ( .A(net_13521), .Z(net_13522) );
CLKBUF_X2 inst_11524 ( .A(net_11371), .Z(net_11372) );
CLKBUF_X2 inst_18989 ( .A(net_18226), .Z(net_18837) );
CLKBUF_X2 inst_18811 ( .A(net_16871), .Z(net_18659) );
INV_X4 inst_5483 ( .ZN(net_733), .A(x2981) );
HA_X1 inst_6694 ( .A(net_3051), .S(net_2871), .CO(net_2870), .B(net_2804) );
NOR2_X2 inst_3373 ( .ZN(net_5552), .A1(net_5336), .A2(net_5334) );
AOI21_X2 inst_8919 ( .B2(net_5843), .ZN(net_5717), .A(net_5715), .B1(net_2729) );
NAND2_X2 inst_4902 ( .ZN(net_3299), .A2(x13330), .A1(x13291) );
CLKBUF_X2 inst_11464 ( .A(net_10198), .Z(net_11312) );
CLKBUF_X2 inst_18072 ( .A(net_17919), .Z(net_17920) );
DFFS_X1 inst_6956 ( .D(net_2511), .CK(net_16329), .SN(x6501), .Q(x926) );
NAND2_X2 inst_4720 ( .A1(net_7373), .ZN(net_1988), .A2(net_1784) );
CLKBUF_X2 inst_16750 ( .A(net_16597), .Z(net_16598) );
CLKBUF_X2 inst_11488 ( .A(net_11335), .Z(net_11336) );
CLKBUF_X2 inst_17699 ( .A(net_17546), .Z(net_17547) );
MUX2_X2 inst_4986 ( .A(net_9028), .Z(net_3966), .B(net_3330), .S(net_622) );
CLKBUF_X2 inst_18980 ( .A(net_18827), .Z(net_18828) );
CLKBUF_X2 inst_18695 ( .A(net_18542), .Z(net_18543) );
INV_X2 inst_6378 ( .ZN(net_1353), .A(net_1352) );
XNOR2_X2 inst_294 ( .A(net_6832), .ZN(net_991), .B(net_990) );
CLKBUF_X2 inst_13510 ( .A(net_13357), .Z(net_13358) );
AOI22_X2 inst_8275 ( .B1(net_8839), .A1(net_8358), .A2(net_6265), .B2(net_6253), .ZN(net_6066) );
AOI22_X2 inst_7842 ( .A2(net_5595), .ZN(net_4667), .B1(net_4666), .B2(net_4388), .A1(net_312) );
CLKBUF_X2 inst_15428 ( .A(net_15275), .Z(net_15276) );
NOR2_X2 inst_3384 ( .ZN(net_5541), .A1(net_5289), .A2(net_5288) );
CLKBUF_X2 inst_11202 ( .A(net_11049), .Z(net_11050) );
SDFF_X2 inst_810 ( .SI(net_8500), .Q(net_8500), .D(net_3958), .SE(net_3884), .CK(net_12252) );
CLKBUF_X2 inst_16540 ( .A(net_10069), .Z(net_16388) );
AOI21_X2 inst_8982 ( .A(net_2146), .ZN(net_2099), .B1(net_1922), .B2(net_1921) );
CLKBUF_X2 inst_16043 ( .A(net_15890), .Z(net_15891) );
CLKBUF_X2 inst_9511 ( .A(net_9358), .Z(net_9359) );
CLKBUF_X2 inst_18895 ( .A(net_18742), .Z(net_18743) );
CLKBUF_X2 inst_9767 ( .A(net_9614), .Z(net_9615) );
OAI21_X2 inst_3035 ( .B2(net_8249), .B1(net_4928), .ZN(net_4843), .A(net_3874) );
CLKBUF_X2 inst_18900 ( .A(net_18747), .Z(net_18748) );
CLKBUF_X2 inst_17694 ( .A(net_17541), .Z(net_17542) );
CLKBUF_X2 inst_14855 ( .A(net_14702), .Z(net_14703) );
CLKBUF_X2 inst_12063 ( .A(net_10218), .Z(net_11911) );
CLKBUF_X2 inst_18015 ( .A(net_17862), .Z(net_17863) );
AOI22_X2 inst_7836 ( .A2(net_5595), .B2(net_4881), .ZN(net_4675), .A1(net_329), .B1(net_247) );
CLKBUF_X2 inst_10010 ( .A(net_9234), .Z(net_9858) );
CLKBUF_X2 inst_14573 ( .A(net_14420), .Z(net_14421) );
CLKBUF_X2 inst_11984 ( .A(net_11831), .Z(net_11832) );
SDFF_X2 inst_481 ( .SI(net_8603), .Q(net_8603), .SE(net_3984), .D(net_3960), .CK(net_13144) );
CLKBUF_X2 inst_16076 ( .A(net_15923), .Z(net_15924) );
INV_X4 inst_5992 ( .A(net_7440), .ZN(net_652) );
CLKBUF_X2 inst_16295 ( .A(net_16142), .Z(net_16143) );
AOI222_X1 inst_8633 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_4363), .B1(net_3987), .C1(net_1329), .A1(x13663) );
CLKBUF_X2 inst_13699 ( .A(net_9405), .Z(net_13547) );
INV_X2 inst_6208 ( .ZN(net_5502), .A(net_5397) );
CLKBUF_X2 inst_16899 ( .A(net_10764), .Z(net_16747) );
CLKBUF_X2 inst_13056 ( .A(net_12903), .Z(net_12904) );
SDFFR_X2 inst_2485 ( .D(net_7366), .SI(net_2555), .SE(net_2288), .QN(net_433), .CK(net_13677), .RN(x6501) );
CLKBUF_X2 inst_16773 ( .A(net_9256), .Z(net_16621) );
AND2_X4 inst_9087 ( .ZN(net_4888), .A2(net_4799), .A1(net_2580) );
CLKBUF_X2 inst_10584 ( .A(net_10431), .Z(net_10432) );
CLKBUF_X2 inst_13353 ( .A(net_9168), .Z(net_13201) );
SDFFR_X2 inst_2217 ( .Q(net_7447), .D(net_7447), .SE(net_2863), .CK(net_12818), .SI(x13605), .RN(x6501) );
CLKBUF_X2 inst_16332 ( .A(net_9712), .Z(net_16180) );
CLKBUF_X2 inst_13707 ( .A(net_13554), .Z(net_13555) );
SDFF_X2 inst_850 ( .SI(net_8663), .Q(net_8663), .D(net_3976), .SE(net_3885), .CK(net_12787) );
CLKBUF_X2 inst_17719 ( .A(net_17566), .Z(net_17567) );
CLKBUF_X2 inst_11175 ( .A(net_9509), .Z(net_11023) );
CLKBUF_X2 inst_12642 ( .A(net_12489), .Z(net_12490) );
CLKBUF_X2 inst_16912 ( .A(net_16759), .Z(net_16760) );
CLKBUF_X2 inst_17444 ( .A(net_17291), .Z(net_17292) );
CLKBUF_X2 inst_14485 ( .A(net_14332), .Z(net_14333) );
SDFFR_X2 inst_2438 ( .D(net_4465), .SE(net_2313), .SI(net_422), .Q(net_422), .CK(net_14815), .RN(x6501) );
CLKBUF_X2 inst_15577 ( .A(net_9093), .Z(net_15425) );
CLKBUF_X2 inst_10391 ( .A(net_9279), .Z(net_10239) );
INV_X4 inst_5479 ( .ZN(net_832), .A(net_740) );
XNOR2_X2 inst_237 ( .ZN(net_1240), .B(net_854), .A(net_532) );
SDFFR_X2 inst_2543 ( .QN(net_6369), .SE(net_2147), .SI(net_1957), .D(net_933), .CK(net_18141), .RN(x6501) );
SDFFR_X1 inst_2772 ( .Q(net_7278), .D(net_2785), .SI(net_1945), .SE(net_1327), .CK(net_14774), .RN(x6501) );
CLKBUF_X2 inst_11449 ( .A(net_9285), .Z(net_11297) );
AOI221_X2 inst_8836 ( .B1(net_8069), .C1(net_7865), .B2(net_6107), .ZN(net_6021), .C2(net_4400), .A(net_4293) );
CLKBUF_X2 inst_17234 ( .A(net_17081), .Z(net_17082) );
CLKBUF_X2 inst_13178 ( .A(net_13025), .Z(net_13026) );
AOI22_X2 inst_8056 ( .A1(net_7968), .B1(net_7798), .A2(net_6092), .B2(net_6091), .ZN(net_4085) );
CLKBUF_X2 inst_17667 ( .A(net_17514), .Z(net_17515) );
XOR2_X2 inst_51 ( .A(net_7572), .B(net_3014), .Z(net_997) );
SDFF_X2 inst_813 ( .SI(net_8503), .Q(net_8503), .D(net_3956), .SE(net_3884), .CK(net_10060) );
CLKBUF_X2 inst_17081 ( .A(net_16928), .Z(net_16929) );
CLKBUF_X2 inst_10379 ( .A(net_10226), .Z(net_10227) );
HA_X1 inst_6691 ( .S(net_2923), .CO(net_2922), .A(net_2921), .B(net_2864) );
CLKBUF_X2 inst_14874 ( .A(net_9952), .Z(net_14722) );
CLKBUF_X2 inst_13373 ( .A(net_13220), .Z(net_13221) );
CLKBUF_X2 inst_11195 ( .A(net_10696), .Z(net_11043) );
SDFF_X2 inst_1837 ( .D(net_7277), .SI(net_6894), .Q(net_6894), .SE(net_6284), .CK(net_17362) );
CLKBUF_X2 inst_18527 ( .A(net_18374), .Z(net_18375) );
CLKBUF_X2 inst_13198 ( .A(net_11132), .Z(net_13046) );
AND2_X4 inst_9100 ( .ZN(net_2543), .A2(net_2268), .A1(net_2261) );
INV_X4 inst_5686 ( .ZN(net_2735), .A(net_161) );
CLKBUF_X2 inst_10944 ( .A(net_10791), .Z(net_10792) );
NOR3_X2 inst_3291 ( .A1(net_2400), .ZN(net_2341), .A3(net_2180), .A2(net_1992) );
XOR2_X2 inst_64 ( .A(net_972), .B(net_945), .Z(net_926) );
CLKBUF_X2 inst_15904 ( .A(net_11902), .Z(net_15752) );
CLKBUF_X2 inst_13964 ( .A(net_11554), .Z(net_13812) );
SDFF_X2 inst_743 ( .Q(net_8808), .D(net_8808), .SI(net_3940), .SE(net_3879), .CK(net_10335) );
SDFFR_X2 inst_2106 ( .SI(net_7406), .Q(net_7406), .SE(net_6198), .D(net_5734), .CK(net_9387), .RN(x6501) );
NAND2_X4 inst_4051 ( .ZN(net_2146), .A2(net_1748), .A1(net_478) );
SDFFR_X1 inst_2723 ( .SI(net_9034), .Q(net_9034), .D(net_7463), .SE(net_3208), .CK(net_10667), .RN(x6501) );
CLKBUF_X2 inst_18825 ( .A(net_16329), .Z(net_18673) );
AND2_X4 inst_9141 ( .A2(net_7482), .A1(net_7480), .ZN(net_1655) );
NAND2_X2 inst_4265 ( .A1(net_6914), .A2(net_5247), .ZN(net_5195) );
AOI222_X1 inst_8628 ( .B2(net_8236), .B1(net_4891), .C2(net_4889), .A1(net_4803), .ZN(net_4796), .C1(net_4459), .A2(net_2873) );
SDFF_X2 inst_1809 ( .D(net_7264), .SI(net_6841), .Q(net_6841), .SE(net_6282), .CK(net_17421) );
HA_X1 inst_6664 ( .A(net_7442), .S(net_3532), .CO(net_3531), .B(net_3232) );
AOI22_X2 inst_8272 ( .B1(net_8691), .A1(net_8654), .B2(net_6109), .A2(net_3857), .ZN(net_3767) );
CLKBUF_X2 inst_14602 ( .A(net_14449), .Z(net_14450) );
CLKBUF_X2 inst_12172 ( .A(net_10679), .Z(net_12020) );
CLKBUF_X2 inst_11866 ( .A(net_11713), .Z(net_11714) );
NAND2_X2 inst_4344 ( .A1(net_7146), .A2(net_5166), .ZN(net_5113) );
AOI22_X2 inst_8111 ( .B1(net_8213), .A1(net_7703), .B2(net_6099), .A2(net_4399), .ZN(net_4036) );
AOI22_X2 inst_8541 ( .B1(net_6726), .A1(net_6693), .B2(net_6202), .A2(net_3520), .ZN(net_3399) );
CLKBUF_X2 inst_15404 ( .A(net_13334), .Z(net_15252) );
CLKBUF_X2 inst_14717 ( .A(net_14564), .Z(net_14565) );
CLKBUF_X2 inst_16794 ( .A(net_16641), .Z(net_16642) );
NAND3_X2 inst_4011 ( .ZN(net_1591), .A1(net_1058), .A3(net_1057), .A2(x12780) );
CLKBUF_X2 inst_17992 ( .A(net_17839), .Z(net_17840) );
CLKBUF_X2 inst_11478 ( .A(net_9383), .Z(net_11326) );
CLKBUF_X2 inst_10432 ( .A(net_10279), .Z(net_10280) );
CLKBUF_X2 inst_15556 ( .A(net_12054), .Z(net_15404) );
CLKBUF_X2 inst_17763 ( .A(net_9428), .Z(net_17611) );
CLKBUF_X2 inst_14609 ( .A(net_14456), .Z(net_14457) );
INV_X2 inst_6445 ( .A(net_6354), .ZN(net_2126) );
CLKBUF_X2 inst_17322 ( .A(net_17169), .Z(net_17170) );
AOI22_X2 inst_8045 ( .A1(net_7967), .B1(net_7797), .A2(net_6092), .B2(net_6091), .ZN(net_4095) );
DFFR_X1 inst_7436 ( .QN(net_8916), .D(net_4848), .CK(net_13978), .RN(x6501) );
CLKBUF_X2 inst_11689 ( .A(net_11536), .Z(net_11537) );
OAI21_X4 inst_2980 ( .B2(net_4926), .ZN(net_3537), .B1(net_3262), .A(net_3189) );
INV_X4 inst_5197 ( .A(net_2527), .ZN(net_2526) );
CLKBUF_X2 inst_18861 ( .A(net_13269), .Z(net_18709) );
CLKBUF_X2 inst_10184 ( .A(net_10031), .Z(net_10032) );
SDFF_X2 inst_915 ( .SI(net_8734), .Q(net_8734), .SE(net_6195), .D(net_3940), .CK(net_13460) );
CLKBUF_X2 inst_9869 ( .A(net_9716), .Z(net_9717) );
NAND2_X2 inst_4416 ( .A1(net_6855), .A2(net_5016), .ZN(net_5011) );
CLKBUF_X2 inst_10008 ( .A(net_9855), .Z(net_9856) );
INV_X4 inst_5660 ( .A(net_7572), .ZN(net_582) );
CLKBUF_X2 inst_16343 ( .A(net_12747), .Z(net_16191) );
CLKBUF_X2 inst_14017 ( .A(net_13864), .Z(net_13865) );
CLKBUF_X2 inst_16096 ( .A(net_11903), .Z(net_15944) );
CLKBUF_X2 inst_9552 ( .A(net_9399), .Z(net_9400) );
CLKBUF_X2 inst_14703 ( .A(net_14550), .Z(net_14551) );
CLKBUF_X2 inst_12591 ( .A(net_12438), .Z(net_12439) );
NAND2_X2 inst_4807 ( .ZN(net_1625), .A2(net_855), .A1(net_839) );
SDFF_X2 inst_1668 ( .SI(net_7766), .Q(net_7766), .D(net_2715), .SE(net_2560), .CK(net_14260) );
CLKBUF_X2 inst_16432 ( .A(net_16279), .Z(net_16280) );
CLKBUF_X2 inst_11169 ( .A(net_9699), .Z(net_11017) );
CLKBUF_X2 inst_9987 ( .A(net_9834), .Z(net_9835) );
CLKBUF_X2 inst_15425 ( .A(net_15272), .Z(net_15273) );
NAND2_X2 inst_4811 ( .ZN(net_2525), .A1(net_1283), .A2(net_806) );
CLKBUF_X2 inst_15935 ( .A(net_11894), .Z(net_15783) );
CLKBUF_X2 inst_11942 ( .A(net_11789), .Z(net_11790) );
DFFR_X2 inst_7068 ( .QN(net_7416), .D(net_4203), .CK(net_12372), .RN(x6501) );
CLKBUF_X2 inst_18726 ( .A(net_18573), .Z(net_18574) );
XNOR2_X2 inst_293 ( .B(net_3194), .ZN(net_998), .A(net_540) );
NAND2_X2 inst_4741 ( .ZN(net_2722), .A2(net_1586), .A1(net_972) );
CLKBUF_X2 inst_11078 ( .A(net_10854), .Z(net_10926) );
NAND4_X2 inst_3744 ( .ZN(net_4286), .A1(net_4052), .A2(net_4051), .A3(net_4050), .A4(net_4049) );
CLKBUF_X2 inst_15346 ( .A(net_9798), .Z(net_15194) );
CLKBUF_X2 inst_17154 ( .A(net_9574), .Z(net_17002) );
INV_X4 inst_5402 ( .ZN(net_2520), .A(net_880) );
CLKBUF_X2 inst_18976 ( .A(net_18823), .Z(net_18824) );
OAI221_X2 inst_2953 ( .C2(net_8234), .B1(net_7577), .B2(net_4971), .ZN(net_4929), .C1(net_4928), .A(net_3112) );
CLKBUF_X2 inst_13000 ( .A(net_12847), .Z(net_12848) );
CLKBUF_X2 inst_17614 ( .A(net_17461), .Z(net_17462) );
AOI22_X2 inst_8219 ( .B1(net_8795), .A1(net_8536), .A2(net_3861), .B2(net_3860), .ZN(net_3817) );
XOR2_X1 inst_98 ( .B(net_1444), .Z(net_1314), .A(net_1078) );
OAI21_X2 inst_3087 ( .ZN(net_3037), .B2(net_2859), .A(net_2025), .B1(net_1835) );
SDFF_X2 inst_959 ( .SI(net_7317), .Q(net_6691), .D(net_6691), .SE(net_3125), .CK(net_9886) );
CLKBUF_X2 inst_10102 ( .A(net_9949), .Z(net_9950) );
CLKBUF_X2 inst_14611 ( .A(net_13948), .Z(net_14459) );
CLKBUF_X2 inst_18397 ( .A(net_18244), .Z(net_18245) );
CLKBUF_X2 inst_13343 ( .A(net_13190), .Z(net_13191) );
SDFF_X2 inst_605 ( .SI(net_8400), .Q(net_8400), .SE(net_3969), .D(net_3952), .CK(net_10360) );
CLKBUF_X2 inst_9998 ( .A(net_9845), .Z(net_9846) );
DFFR_X1 inst_7481 ( .QN(net_7427), .D(net_4211), .CK(net_12385), .RN(x6501) );
OR3_X4 inst_2799 ( .ZN(net_2943), .A1(net_2425), .A3(net_2308), .A2(net_1819) );
CLKBUF_X2 inst_10988 ( .A(net_9446), .Z(net_10836) );
SDFF_X2 inst_2048 ( .SI(net_7908), .Q(net_7908), .D(net_2721), .SE(net_2461), .CK(net_15805) );
OAI222_X2 inst_2948 ( .ZN(net_3890), .A2(net_3889), .B2(net_3888), .C2(net_3887), .A1(net_2175), .B1(net_1665), .C1(net_657) );
AOI22_X2 inst_7900 ( .ZN(net_4529), .B1(net_4528), .A2(net_4515), .B2(net_4388), .A1(net_2800) );
CLKBUF_X2 inst_10396 ( .A(net_9829), .Z(net_10244) );
CLKBUF_X2 inst_11643 ( .A(net_11234), .Z(net_11491) );
CLKBUF_X2 inst_13850 ( .A(net_13697), .Z(net_13698) );
SDFF_X2 inst_1931 ( .SI(net_8060), .Q(net_8060), .D(net_2575), .SE(net_2508), .CK(net_15958) );
NAND2_X2 inst_4735 ( .ZN(net_2702), .A2(net_1586), .A1(net_931) );
INV_X16 inst_6631 ( .ZN(net_3864), .A(net_3372) );
CLKBUF_X2 inst_11926 ( .A(net_11773), .Z(net_11774) );
AOI22_X2 inst_8402 ( .A1(net_8600), .B1(net_8415), .A2(net_3864), .B2(net_3863), .ZN(net_3650) );
OAI21_X2 inst_3002 ( .B2(net_5902), .ZN(net_5891), .A(net_5823), .B1(net_728) );
CLKBUF_X2 inst_13007 ( .A(net_11622), .Z(net_12855) );
NAND2_X2 inst_4389 ( .A1(net_7123), .A2(net_5166), .ZN(net_5068) );
DFF_X1 inst_6828 ( .Q(net_6448), .D(net_3620), .CK(net_17914) );
CLKBUF_X2 inst_15153 ( .A(net_15000), .Z(net_15001) );
OAI22_X2 inst_2940 ( .B2(net_2147), .ZN(net_1997), .A1(net_1996), .A2(net_1710), .B1(net_688) );
CLKBUF_X2 inst_16391 ( .A(net_16238), .Z(net_16239) );
CLKBUF_X2 inst_11855 ( .A(net_11702), .Z(net_11703) );
DFFR_X1 inst_7533 ( .D(net_918), .Q(net_397), .CK(net_18734), .RN(x6501) );
CLKBUF_X2 inst_9383 ( .A(net_9157), .Z(net_9231) );
INV_X2 inst_6606 ( .A(net_6169), .ZN(net_6165) );
CLKBUF_X2 inst_11267 ( .A(net_11114), .Z(net_11115) );
CLKBUF_X2 inst_15048 ( .A(net_9130), .Z(net_14896) );
DFFR_X2 inst_7022 ( .QN(net_6291), .D(net_5707), .CK(net_13869), .RN(x6501) );
NOR2_X2 inst_3474 ( .ZN(net_5031), .A2(net_5027), .A1(net_1139) );
CLKBUF_X2 inst_16136 ( .A(net_15983), .Z(net_15984) );
CLKBUF_X2 inst_12328 ( .A(net_12175), .Z(net_12176) );
SDFF_X2 inst_578 ( .Q(net_8844), .D(net_8844), .SE(net_3964), .SI(net_3952), .CK(net_10363) );
CLKBUF_X2 inst_17251 ( .A(net_17098), .Z(net_17099) );
CLKBUF_X2 inst_17913 ( .A(net_17760), .Z(net_17761) );
CLKBUF_X2 inst_16129 ( .A(net_15976), .Z(net_15977) );
CLKBUF_X2 inst_14197 ( .A(net_14044), .Z(net_14045) );
CLKBUF_X2 inst_13063 ( .A(net_12910), .Z(net_12911) );
CLKBUF_X2 inst_17873 ( .A(net_17720), .Z(net_17721) );
CLKBUF_X2 inst_15164 ( .A(net_13150), .Z(net_15012) );
DFFR_X2 inst_7317 ( .D(net_6827), .QN(net_6824), .CK(net_15092), .RN(x6501) );
CLKBUF_X2 inst_18355 ( .A(net_18202), .Z(net_18203) );
SDFF_X2 inst_1498 ( .SI(net_7855), .Q(net_7855), .D(net_2576), .SE(net_2558), .CK(net_16061) );
SDFF_X2 inst_1358 ( .SI(net_7712), .Q(net_7712), .D(net_2702), .SE(net_2559), .CK(net_18870) );
AOI22_X2 inst_8343 ( .B1(net_8811), .A1(net_8552), .A2(net_3861), .B2(net_3860), .ZN(net_3704) );
CLKBUF_X2 inst_17853 ( .A(net_17700), .Z(net_17701) );
CLKBUF_X2 inst_18935 ( .A(net_17951), .Z(net_18783) );
CLKBUF_X2 inst_12456 ( .A(net_12254), .Z(net_12304) );
NAND2_X2 inst_4775 ( .A2(net_2528), .ZN(net_1799), .A1(net_1618) );
CLKBUF_X2 inst_16303 ( .A(net_16150), .Z(net_16151) );
CLKBUF_X2 inst_10831 ( .A(net_10678), .Z(net_10679) );
NAND2_X2 inst_4450 ( .ZN(net_4977), .A2(net_4795), .A1(net_4529) );
CLKBUF_X2 inst_12817 ( .A(net_11489), .Z(net_12665) );
CLKBUF_X2 inst_17856 ( .A(net_17703), .Z(net_17704) );
CLKBUF_X2 inst_12460 ( .A(net_12307), .Z(net_12308) );
OAI211_X2 inst_3182 ( .C2(net_8237), .ZN(net_5587), .A(net_5455), .C1(net_4954), .B(net_4677) );
CLKBUF_X2 inst_14557 ( .A(net_14404), .Z(net_14405) );
OR2_X2 inst_2866 ( .ZN(net_5921), .A2(net_5920), .A1(net_2412) );
DFF_X1 inst_6805 ( .Q(net_8222), .D(net_4423), .CK(net_16561) );
CLKBUF_X2 inst_11528 ( .A(net_9415), .Z(net_11376) );
CLKBUF_X2 inst_11546 ( .A(net_9712), .Z(net_11394) );
INV_X4 inst_5379 ( .ZN(net_1976), .A(net_716) );
SDFF_X2 inst_838 ( .SI(net_8649), .Q(net_8649), .D(net_3974), .SE(net_3885), .CK(net_10140) );
CLKBUF_X2 inst_12905 ( .A(net_11177), .Z(net_12753) );
SDFF_X2 inst_1405 ( .SI(net_7289), .Q(net_7066), .D(net_7066), .SE(net_6280), .CK(net_18402) );
DFF_X1 inst_6811 ( .Q(net_8252), .D(net_4427), .CK(net_17593) );
NAND2_X2 inst_4058 ( .ZN(net_5906), .A2(net_5836), .A1(net_3115) );
DFF_X1 inst_6786 ( .Q(net_7535), .D(net_4584), .CK(net_11957) );
AND2_X2 inst_9172 ( .ZN(net_2751), .A1(net_2493), .A2(net_2382) );
SDFFR_X1 inst_2749 ( .SI(net_9033), .Q(net_9033), .D(net_7462), .SE(net_3208), .CK(net_10641), .RN(x6501) );
INV_X4 inst_5584 ( .A(net_7386), .ZN(net_596) );
DFFS_X1 inst_6963 ( .Q(net_8263), .D(net_959), .CK(net_18486), .SN(x6501) );
CLKBUF_X2 inst_19065 ( .A(net_18912), .Z(net_18913) );
AOI221_X2 inst_8823 ( .B1(net_8044), .C1(net_7840), .B2(net_6107), .ZN(net_5995), .C2(net_4400), .A(net_4310) );
CLKBUF_X2 inst_11118 ( .A(net_10965), .Z(net_10966) );
CLKBUF_X2 inst_14647 ( .A(net_14494), .Z(net_14495) );
INV_X4 inst_5567 ( .A(net_7510), .ZN(net_3388) );
SDFF_X2 inst_2013 ( .SI(net_7909), .Q(net_7909), .D(net_2585), .SE(net_2461), .CK(net_15808) );
NAND2_X2 inst_4506 ( .A2(net_6800), .A1(net_6272), .ZN(net_4359) );
SDFFR_X1 inst_2756 ( .QN(net_7581), .D(net_3957), .SE(net_3144), .SI(net_755), .CK(net_10959), .RN(x6501) );
CLKBUF_X2 inst_10071 ( .A(net_9918), .Z(net_9919) );
SDFF_X2 inst_492 ( .SI(net_8616), .Q(net_8616), .SE(net_3984), .D(net_3942), .CK(net_12630) );
AOI222_X1 inst_8635 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_4229), .B1(net_3583), .C1(net_3581), .A1(x13742) );
DFFR_X2 inst_7229 ( .QN(net_8215), .D(net_2254), .CK(net_17307), .RN(x6501) );
INV_X4 inst_5414 ( .ZN(net_866), .A(net_865) );
CLKBUF_X2 inst_18298 ( .A(net_18145), .Z(net_18146) );
CLKBUF_X2 inst_12589 ( .A(net_12436), .Z(net_12437) );
CLKBUF_X2 inst_12292 ( .A(net_12139), .Z(net_12140) );
XOR2_X1 inst_82 ( .Z(net_3049), .B(net_3048), .A(net_2922) );
NAND2_X2 inst_4335 ( .A1(net_7143), .A2(net_5166), .ZN(net_5122) );
NAND2_X2 inst_4187 ( .ZN(net_5314), .A1(net_5185), .A2(net_4985) );
NAND2_X2 inst_4239 ( .A1(net_6902), .A2(net_5247), .ZN(net_5221) );
CLKBUF_X2 inst_15586 ( .A(net_15433), .Z(net_15434) );
DFFR_X2 inst_7335 ( .Q(net_7319), .CK(net_11364), .D(x13100), .RN(x6501) );
CLKBUF_X2 inst_12171 ( .A(net_12018), .Z(net_12019) );
SDFF_X2 inst_1121 ( .D(net_7326), .SI(net_6568), .Q(net_6568), .SE(net_3070), .CK(net_11316) );
CLKBUF_X2 inst_12185 ( .A(net_12032), .Z(net_12033) );
AOI21_X2 inst_8932 ( .B2(net_5843), .ZN(net_5678), .A(net_5677), .B1(x324) );
OAI211_X2 inst_3187 ( .ZN(net_4927), .B(net_4926), .C1(net_4922), .A(net_4837), .C2(net_4836) );
CLKBUF_X2 inst_18213 ( .A(net_18060), .Z(net_18061) );
CLKBUF_X2 inst_11053 ( .A(net_10900), .Z(net_10901) );
CLKBUF_X2 inst_17294 ( .A(net_17141), .Z(net_17142) );
XNOR2_X2 inst_307 ( .A(net_1864), .ZN(net_965), .B(net_203) );
AOI22_X2 inst_8411 ( .A1(net_8602), .B1(net_8417), .A2(net_3864), .B2(net_3863), .ZN(net_3641) );
AOI22_X2 inst_8292 ( .A1(net_8620), .B1(net_8435), .A2(net_3864), .B2(net_3863), .ZN(net_3750) );
CLKBUF_X2 inst_12663 ( .A(net_9559), .Z(net_12511) );
CLKBUF_X2 inst_18291 ( .A(net_16117), .Z(net_18139) );
SDFF_X2 inst_2034 ( .SI(net_7786), .Q(net_7786), .D(net_2589), .SE(net_2459), .CK(net_18341) );
CLKBUF_X2 inst_16354 ( .A(net_12756), .Z(net_16202) );
SDFF_X2 inst_717 ( .SI(net_8648), .Q(net_8648), .D(net_3958), .SE(net_3885), .CK(net_10993) );
SDFF_X2 inst_1505 ( .SI(net_7865), .Q(net_7865), .D(net_2711), .SE(net_2558), .CK(net_14286) );
CLKBUF_X2 inst_15097 ( .A(net_14944), .Z(net_14945) );
CLKBUF_X2 inst_10439 ( .A(net_10286), .Z(net_10287) );
AOI22_X2 inst_8460 ( .B1(net_6539), .A1(net_6506), .A2(net_6137), .B2(net_6104), .ZN(net_3480) );
CLKBUF_X2 inst_11557 ( .A(net_11404), .Z(net_11405) );
DFFR_X2 inst_7166 ( .QN(net_8944), .D(net_2647), .CK(net_16308), .RN(x6501) );
CLKBUF_X2 inst_19037 ( .A(net_18884), .Z(net_18885) );
CLKBUF_X2 inst_16693 ( .A(net_16540), .Z(net_16541) );
AOI22_X2 inst_7944 ( .B1(net_8191), .A1(net_7681), .B2(net_6099), .A2(net_4399), .ZN(net_4181) );
NAND4_X2 inst_3686 ( .ZN(net_4451), .A4(net_4351), .A1(net_3851), .A2(net_3850), .A3(net_3849) );
CLKBUF_X2 inst_15956 ( .A(net_15803), .Z(net_15804) );
NAND4_X2 inst_3842 ( .ZN(net_1841), .A1(net_1558), .A4(net_1555), .A2(net_1220), .A3(net_998) );
CLKBUF_X2 inst_12186 ( .A(net_10260), .Z(net_12034) );
SDFF_X2 inst_1703 ( .SI(net_7705), .Q(net_7705), .D(net_2585), .SE(net_2559), .CK(net_18522) );
INV_X4 inst_5886 ( .A(net_9009), .ZN(net_915) );
INV_X2 inst_6566 ( .A(net_6329), .ZN(net_489) );
DFFR_X2 inst_7167 ( .QN(net_8943), .D(net_2648), .CK(net_16304), .RN(x6501) );
CLKBUF_X2 inst_18122 ( .A(net_17969), .Z(net_17970) );
CLKBUF_X2 inst_14894 ( .A(net_9960), .Z(net_14742) );
CLKBUF_X2 inst_14139 ( .A(net_13986), .Z(net_13987) );
CLKBUF_X2 inst_13680 ( .A(net_12593), .Z(net_13528) );
AOI22_X2 inst_7788 ( .A2(net_6187), .B2(net_5535), .ZN(net_4812), .B1(net_467), .A1(net_198) );
CLKBUF_X2 inst_16358 ( .A(net_16205), .Z(net_16206) );
AOI21_X2 inst_8934 ( .B2(net_5784), .ZN(net_5672), .A(net_5671), .B1(x534) );
SDFF_X2 inst_614 ( .SI(net_8377), .Q(net_8377), .SE(net_3969), .D(net_3947), .CK(net_12448) );
AND2_X4 inst_9080 ( .ZN(net_3125), .A2(net_2940), .A1(net_2901) );
CLKBUF_X2 inst_12197 ( .A(net_12044), .Z(net_12045) );
SDFF_X2 inst_1896 ( .D(net_7286), .SI(net_7023), .Q(net_7023), .SE(net_6277), .CK(net_16182) );
SDFF_X2 inst_1031 ( .SI(net_7312), .Q(net_6719), .D(net_6719), .SE(net_3124), .CK(net_9865) );
SDFF_X2 inst_945 ( .SI(net_7327), .Q(net_6701), .D(net_6701), .SE(net_3125), .CK(net_9107) );
CLKBUF_X2 inst_17012 ( .A(net_16859), .Z(net_16860) );
SDFF_X2 inst_369 ( .SI(net_8320), .Q(net_8320), .SE(net_3978), .D(net_3942), .CK(net_12803) );
SDFF_X2 inst_1900 ( .D(net_7292), .SI(net_7029), .Q(net_7029), .SE(net_6277), .CK(net_14874) );
CLKBUF_X2 inst_15044 ( .A(net_9590), .Z(net_14892) );
CLKBUF_X2 inst_12899 ( .A(net_9078), .Z(net_12747) );
CLKBUF_X2 inst_12850 ( .A(net_12697), .Z(net_12698) );
INV_X4 inst_5695 ( .ZN(net_723), .A(net_342) );
OAI22_X2 inst_2916 ( .ZN(net_3540), .A2(net_3538), .B2(net_3537), .A1(net_1623), .B1(net_1476) );
SDFF_X2 inst_1286 ( .Q(net_7829), .D(net_7829), .SI(net_2749), .SE(net_2730), .CK(net_16516) );
AOI221_X2 inst_8812 ( .C2(net_5609), .B2(net_5520), .A(net_4834), .ZN(net_4716), .C1(net_358), .B1(net_288) );
CLKBUF_X2 inst_18599 ( .A(net_14921), .Z(net_18447) );
XOR2_X1 inst_77 ( .Z(net_3275), .B(net_3274), .A(net_3168) );
INV_X2 inst_6399 ( .ZN(net_1159), .A(net_1158) );
AOI22_X2 inst_8224 ( .B1(net_8574), .A1(net_8463), .A2(net_6263), .B2(net_6262), .ZN(net_3813) );
CLKBUF_X2 inst_17010 ( .A(net_16857), .Z(net_16858) );
CLKBUF_X2 inst_17435 ( .A(net_17282), .Z(net_17283) );
CLKBUF_X2 inst_13328 ( .A(net_13175), .Z(net_13176) );
CLKBUF_X2 inst_11710 ( .A(net_9593), .Z(net_11558) );
DFFR_X2 inst_7086 ( .QN(net_7652), .D(net_3890), .CK(net_12675), .RN(x6501) );
CLKBUF_X2 inst_9642 ( .A(net_9489), .Z(net_9490) );
CLKBUF_X2 inst_18483 ( .A(net_18330), .Z(net_18331) );
CLKBUF_X2 inst_15713 ( .A(net_10117), .Z(net_15561) );
CLKBUF_X2 inst_11881 ( .A(net_11728), .Z(net_11729) );
CLKBUF_X2 inst_19070 ( .A(net_18917), .Z(net_18918) );
CLKBUF_X2 inst_13553 ( .A(net_13400), .Z(net_13401) );
CLKBUF_X2 inst_14691 ( .A(net_14538), .Z(net_14539) );
CLKBUF_X2 inst_9637 ( .A(net_9284), .Z(net_9485) );
CLKBUF_X2 inst_19199 ( .A(net_19046), .Z(net_19047) );
SDFF_X2 inst_1234 ( .Q(net_7837), .D(net_7837), .SE(net_2730), .SI(net_2716), .CK(net_17106) );
CLKBUF_X2 inst_10040 ( .A(net_9887), .Z(net_9888) );
CLKBUF_X2 inst_16564 ( .A(net_16411), .Z(net_16412) );
SDFFR_X2 inst_2398 ( .SI(net_7376), .SE(net_2723), .D(net_2352), .QN(net_157), .CK(net_15037), .RN(x6501) );
SDFFR_X2 inst_2595 ( .D(net_7379), .QN(net_7239), .SI(net_1941), .SE(net_1379), .CK(net_14738), .RN(x6501) );
INV_X4 inst_5614 ( .A(net_7493), .ZN(net_4714) );
CLKBUF_X2 inst_11938 ( .A(net_10300), .Z(net_11786) );
CLKBUF_X2 inst_9400 ( .A(net_9149), .Z(net_9248) );
SDFFR_X2 inst_2371 ( .SI(net_5943), .SE(net_2260), .Q(net_350), .D(net_350), .CK(net_11571), .RN(x6501) );
OAI22_X2 inst_2939 ( .A2(net_2250), .ZN(net_2006), .A1(net_1291), .B1(net_1290), .B2(net_1155) );
DFF_X1 inst_6818 ( .QN(net_8233), .D(net_4448), .CK(net_14458) );
SDFF_X2 inst_1223 ( .Q(net_7959), .D(net_7959), .SE(net_2755), .SI(net_2719), .CK(net_18822) );
SDFFR_X1 inst_2785 ( .D(net_7377), .Q(net_7274), .SI(net_1952), .SE(net_1327), .CK(net_17413), .RN(x6501) );
CLKBUF_X2 inst_13636 ( .A(net_13405), .Z(net_13484) );
INV_X2 inst_6574 ( .ZN(net_795), .A(net_222) );
CLKBUF_X2 inst_18578 ( .A(net_18425), .Z(net_18426) );
SDFF_X2 inst_681 ( .Q(net_8688), .D(net_8688), .SI(net_3956), .SE(net_3935), .CK(net_10914) );
INV_X4 inst_5432 ( .ZN(net_1146), .A(net_831) );
CLKBUF_X2 inst_13785 ( .A(net_13632), .Z(net_13633) );
NAND2_X2 inst_4886 ( .A2(net_7378), .ZN(net_711), .A1(net_167) );
CLKBUF_X2 inst_15376 ( .A(net_14077), .Z(net_15224) );
SDFF_X2 inst_2010 ( .SI(net_7778), .Q(net_7778), .D(net_2708), .SE(net_2459), .CK(net_15477) );
CLKBUF_X2 inst_13181 ( .A(net_13028), .Z(net_13029) );
CLKBUF_X2 inst_15604 ( .A(net_15451), .Z(net_15452) );
CLKBUF_X2 inst_11575 ( .A(net_11422), .Z(net_11423) );
INV_X4 inst_5547 ( .A(net_1266), .ZN(net_1091) );
SDFF_X2 inst_871 ( .Q(net_8581), .D(net_8581), .SI(net_3954), .SE(net_3878), .CK(net_10054) );
SDFFR_X1 inst_2684 ( .SI(net_7545), .SE(net_5043), .CK(net_9687), .RN(x6501), .Q(x3996), .D(x3996) );
INV_X2 inst_6320 ( .ZN(net_3343), .A(net_3288) );
DFF_X1 inst_6842 ( .Q(net_6432), .D(net_3605), .CK(net_17971) );
SDFF_X2 inst_1171 ( .D(net_7330), .SI(net_6506), .Q(net_6506), .SE(net_3071), .CK(net_11306) );
CLKBUF_X2 inst_18770 ( .A(net_18617), .Z(net_18618) );
INV_X4 inst_5274 ( .ZN(net_1963), .A(net_1452) );
INV_X4 inst_5493 ( .ZN(net_720), .A(net_719) );
INV_X4 inst_5616 ( .A(net_6382), .ZN(net_1489) );
AOI22_X2 inst_8192 ( .B1(net_8754), .A1(net_8384), .A2(net_3867), .B2(net_3866), .ZN(net_3842) );
INV_X4 inst_5766 ( .A(net_7504), .ZN(net_3236) );
CLKBUF_X2 inst_18026 ( .A(net_17873), .Z(net_17874) );
SDFFR_X2 inst_2594 ( .D(net_7384), .QN(net_7244), .SI(net_1942), .SE(net_1379), .CK(net_14741), .RN(x6501) );
INV_X4 inst_5113 ( .ZN(net_5775), .A(net_4704) );
CLKBUF_X2 inst_16474 ( .A(net_16321), .Z(net_16322) );
CLKBUF_X2 inst_14052 ( .A(net_13899), .Z(net_13900) );
NAND3_X2 inst_3976 ( .ZN(net_2096), .A3(net_1816), .A2(net_1525), .A1(net_1288) );
CLKBUF_X2 inst_11773 ( .A(net_11620), .Z(net_11621) );
CLKBUF_X2 inst_9444 ( .A(net_9116), .Z(net_9292) );
SDFF_X2 inst_1119 ( .D(net_7323), .SI(net_6565), .Q(net_6565), .SE(net_3070), .CK(net_11345) );
CLKBUF_X2 inst_15430 ( .A(net_14723), .Z(net_15278) );
CLKBUF_X2 inst_14748 ( .A(net_9224), .Z(net_14596) );
NAND4_X2 inst_3699 ( .A4(net_6226), .A1(net_6225), .ZN(net_4438), .A2(net_3768), .A3(net_3767) );
INV_X4 inst_5082 ( .ZN(net_5744), .A(net_5717) );
CLKBUF_X2 inst_9684 ( .A(net_9531), .Z(net_9532) );
INV_X8 inst_5050 ( .A(net_6194), .ZN(net_6193) );
CLKBUF_X2 inst_10947 ( .A(net_10794), .Z(net_10795) );
CLKBUF_X2 inst_17310 ( .A(net_17157), .Z(net_17158) );
AND2_X4 inst_9112 ( .ZN(net_1935), .A1(net_1750), .A2(net_1749) );
MUX2_X2 inst_4925 ( .Z(net_3554), .S(net_3552), .B(net_1243), .A(net_956) );
DFFR_X2 inst_7021 ( .QN(net_6307), .D(net_5710), .CK(net_16934), .RN(x6501) );
NAND2_X2 inst_4457 ( .ZN(net_4948), .A2(net_4835), .A1(net_4507) );
INV_X4 inst_6133 ( .A(net_7430), .ZN(net_3098) );
SDFF_X2 inst_903 ( .SI(net_8720), .Q(net_8720), .SE(net_6195), .D(net_3944), .CK(net_10816) );
CLKBUF_X2 inst_14806 ( .A(net_14653), .Z(net_14654) );
SDFF_X2 inst_1725 ( .Q(net_7996), .D(net_7996), .SI(net_2718), .SE(net_2542), .CK(net_15579) );
INV_X4 inst_5391 ( .ZN(net_1608), .A(net_1086) );
DFFR_X2 inst_7238 ( .Q(net_7165), .D(net_2190), .CK(net_18719), .RN(x6501) );
AOI222_X1 inst_8607 ( .B2(net_6785), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5816), .A1(net_3173), .C1(x2308) );
AOI222_X1 inst_8602 ( .B2(net_6764), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5822), .A1(net_2564), .C1(x3288) );
CLKBUF_X2 inst_9700 ( .A(net_9547), .Z(net_9548) );
NOR2_X2 inst_3504 ( .ZN(net_2164), .A2(net_1876), .A1(net_1773) );
NAND3_X2 inst_3924 ( .ZN(net_5614), .A1(net_5543), .A3(net_5477), .A2(net_5295) );
CLKBUF_X2 inst_17365 ( .A(net_17212), .Z(net_17213) );
CLKBUF_X2 inst_14408 ( .A(net_14255), .Z(net_14256) );
NAND2_X2 inst_4510 ( .A1(net_6327), .A2(net_6210), .ZN(net_4354) );
CLKBUF_X2 inst_9548 ( .A(net_9395), .Z(net_9396) );
NAND2_X2 inst_4572 ( .ZN(net_3030), .A1(net_3029), .A2(net_3028) );
INV_X4 inst_5189 ( .ZN(net_2743), .A(net_2557) );
CLKBUF_X2 inst_13053 ( .A(net_11019), .Z(net_12901) );
CLKBUF_X2 inst_17995 ( .A(net_17842), .Z(net_17843) );
CLKBUF_X2 inst_17904 ( .A(net_16671), .Z(net_17752) );
CLKBUF_X2 inst_11203 ( .A(net_11050), .Z(net_11051) );
NOR2_X2 inst_3464 ( .A1(net_2768), .ZN(net_2519), .A2(net_2416) );
SDFF_X2 inst_1044 ( .SI(net_7319), .Q(net_6660), .D(net_6660), .SE(net_3126), .CK(net_12016) );
CLKBUF_X2 inst_9233 ( .A(net_9080), .Z(net_9081) );
INV_X2 inst_6187 ( .ZN(net_5798), .A(net_5763) );
CLKBUF_X2 inst_18907 ( .A(net_18754), .Z(net_18755) );
CLKBUF_X2 inst_10309 ( .A(net_10156), .Z(net_10157) );
DFFR_X1 inst_7554 ( .D(net_2731), .Q(net_291), .CK(net_11184), .RN(x6501) );
CLKBUF_X2 inst_9509 ( .A(net_9348), .Z(net_9357) );
CLKBUF_X2 inst_16377 ( .A(net_16224), .Z(net_16225) );
CLKBUF_X2 inst_16086 ( .A(net_13346), .Z(net_15934) );
CLKBUF_X2 inst_14389 ( .A(net_14236), .Z(net_14237) );
CLKBUF_X2 inst_17191 ( .A(net_16473), .Z(net_17039) );
AOI22_X2 inst_8327 ( .A1(net_8624), .B1(net_8439), .A2(net_3864), .B2(net_3863), .ZN(net_3719) );
OAI21_X2 inst_3014 ( .B1(net_7346), .ZN(net_5462), .A(net_5461), .B2(x1130) );
CLKBUF_X2 inst_16396 ( .A(net_16243), .Z(net_16244) );
CLKBUF_X2 inst_15112 ( .A(net_14959), .Z(net_14960) );
INV_X2 inst_6256 ( .A(net_4901), .ZN(net_4723) );
XNOR2_X2 inst_227 ( .A(net_6204), .ZN(net_1359), .B(net_709) );
SDFF_X2 inst_1532 ( .Q(net_7880), .D(net_7880), .SI(net_2708), .SE(net_2543), .CK(net_18275) );
NAND2_X2 inst_4303 ( .A1(net_7093), .A2(net_5164), .ZN(net_5154) );
INV_X4 inst_5861 ( .A(net_8909), .ZN(net_4528) );
SDFFR_X2 inst_2136 ( .SI(net_7197), .Q(net_7197), .D(net_6448), .SE(net_4362), .CK(net_14561), .RN(x6501) );
CLKBUF_X2 inst_16872 ( .A(net_16719), .Z(net_16720) );
OR2_X2 inst_2891 ( .ZN(net_1755), .A2(net_1574), .A1(net_1170) );
CLKBUF_X2 inst_17830 ( .A(net_17677), .Z(net_17678) );
CLKBUF_X2 inst_18491 ( .A(net_17158), .Z(net_18339) );
CLKBUF_X2 inst_17260 ( .A(net_17107), .Z(net_17108) );
DFFR_X1 inst_7557 ( .D(net_384), .QN(net_383), .CK(net_15214), .RN(x6501) );
AOI222_X1 inst_8642 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3931), .B1(net_3226), .C1(net_3224), .A1(x13684) );
INV_X4 inst_6036 ( .A(net_7211), .ZN(net_502) );
CLKBUF_X2 inst_18381 ( .A(net_18228), .Z(net_18229) );
CLKBUF_X2 inst_9944 ( .A(net_9791), .Z(net_9792) );
CLKBUF_X2 inst_17539 ( .A(net_17386), .Z(net_17387) );
INV_X8 inst_5029 ( .ZN(net_3885), .A(net_3302) );
CLKBUF_X2 inst_10200 ( .A(net_9078), .Z(net_10048) );
CLKBUF_X2 inst_18637 ( .A(net_15140), .Z(net_18485) );
CLKBUF_X2 inst_15457 ( .A(net_15304), .Z(net_15305) );
SDFF_X2 inst_581 ( .Q(net_8847), .D(net_8847), .SE(net_3964), .SI(net_3950), .CK(net_10556) );
SDFFR_X2 inst_2551 ( .SI(net_6830), .Q(net_6830), .SE(net_2146), .D(net_681), .CK(net_18693), .RN(x6501) );
XOR2_X2 inst_28 ( .A(net_2104), .Z(net_1224), .B(net_1221) );
NAND2_X2 inst_4407 ( .A1(net_7129), .A2(net_5166), .ZN(net_5050) );
CLKBUF_X2 inst_17928 ( .A(net_10097), .Z(net_17776) );
CLKBUF_X2 inst_16517 ( .A(net_16364), .Z(net_16365) );
CLKBUF_X2 inst_9410 ( .A(net_9161), .Z(net_9258) );
CLKBUF_X2 inst_12656 ( .A(net_10565), .Z(net_12504) );
CLKBUF_X2 inst_9434 ( .A(net_9281), .Z(net_9282) );
CLKBUF_X2 inst_9401 ( .A(net_9248), .Z(net_9249) );
DFFR_X1 inst_7440 ( .QN(net_8928), .D(net_4755), .CK(net_13975), .RN(x6501) );
CLKBUF_X2 inst_15869 ( .A(net_15716), .Z(net_15717) );
SDFF_X2 inst_592 ( .SI(net_8383), .Q(net_8383), .SE(net_3969), .D(net_3945), .CK(net_13049) );
DFFR_X2 inst_7289 ( .Q(net_7302), .D(net_1327), .CK(net_18257), .RN(x6501) );
CLKBUF_X2 inst_13841 ( .A(net_13688), .Z(net_13689) );
INV_X4 inst_5143 ( .ZN(net_3552), .A(net_3277) );
CLKBUF_X2 inst_15118 ( .A(net_14965), .Z(net_14966) );
CLKBUF_X2 inst_16621 ( .A(net_14102), .Z(net_16469) );
CLKBUF_X2 inst_13504 ( .A(net_12006), .Z(net_13352) );
AOI22_X2 inst_7858 ( .A2(net_5260), .ZN(net_4649), .B2(net_4647), .B1(net_2965), .A1(net_2539) );
CLKBUF_X2 inst_14755 ( .A(net_14602), .Z(net_14603) );
CLKBUF_X2 inst_12876 ( .A(net_12723), .Z(net_12724) );
INV_X4 inst_5096 ( .ZN(net_5697), .A(net_5672) );
NAND3_X2 inst_3948 ( .A3(net_6208), .ZN(net_4512), .A2(net_4323), .A1(net_1504) );
CLKBUF_X2 inst_11413 ( .A(net_11260), .Z(net_11261) );
INV_X4 inst_5227 ( .ZN(net_2259), .A(net_2191) );
CLKBUF_X2 inst_16278 ( .A(net_14099), .Z(net_16126) );
CLKBUF_X2 inst_14157 ( .A(net_11025), .Z(net_14005) );
CLKBUF_X2 inst_11808 ( .A(net_11655), .Z(net_11656) );
CLKBUF_X2 inst_18743 ( .A(net_14842), .Z(net_18591) );
SDFF_X2 inst_1301 ( .Q(net_8095), .D(net_8095), .SI(net_2719), .SE(net_2707), .CK(net_18808) );
CLKBUF_X2 inst_14109 ( .A(net_13956), .Z(net_13957) );
SDFF_X2 inst_647 ( .Q(net_8418), .D(net_8418), .SI(net_3960), .SE(net_3934), .CK(net_13113) );
OR2_X4 inst_2830 ( .ZN(net_3311), .A2(net_3219), .A1(net_3019) );
CLKBUF_X2 inst_12871 ( .A(net_10634), .Z(net_12719) );
CLKBUF_X2 inst_18736 ( .A(net_16761), .Z(net_18584) );
INV_X4 inst_5137 ( .ZN(net_3561), .A(net_3526) );
OAI21_X2 inst_2985 ( .ZN(net_5917), .B2(net_5912), .A(net_5803), .B1(net_645) );
CLKBUF_X2 inst_9821 ( .A(net_9668), .Z(net_9669) );
AOI22_X2 inst_8156 ( .B1(net_8053), .A1(net_7849), .B2(net_6107), .A2(net_4400), .ZN(net_3996) );
SDFF_X2 inst_833 ( .SI(net_8642), .Q(net_8642), .D(net_3945), .SE(net_3885), .CK(net_13330) );
CLKBUF_X2 inst_11968 ( .A(net_11815), .Z(net_11816) );
XNOR2_X2 inst_118 ( .ZN(net_3006), .A(net_2858), .B(net_797) );
MUX2_X2 inst_4924 ( .Z(net_4268), .S(net_3875), .A(net_3535), .B(net_3352) );
CLKBUF_X2 inst_12709 ( .A(net_12556), .Z(net_12557) );
CLKBUF_X2 inst_14433 ( .A(net_14280), .Z(net_14281) );
CLKBUF_X2 inst_10781 ( .A(net_10628), .Z(net_10629) );
INV_X2 inst_6591 ( .A(net_6122), .ZN(net_6121) );
SDFF_X2 inst_2037 ( .SI(net_7772), .Q(net_7772), .D(net_2721), .SE(net_2459), .CK(net_15729) );
AOI22_X2 inst_8578 ( .B1(net_2666), .A2(net_1588), .ZN(net_1519), .A1(net_1518), .B2(net_1517) );
CLKBUF_X2 inst_13532 ( .A(net_9618), .Z(net_13380) );
DFFS_X1 inst_6930 ( .D(net_6145), .CK(net_16359), .SN(x6501), .Q(x856) );
AND2_X4 inst_9102 ( .ZN(net_2381), .A2(net_2188), .A1(net_1175) );
CLKBUF_X2 inst_15343 ( .A(net_13372), .Z(net_15191) );
CLKBUF_X2 inst_12276 ( .A(net_12123), .Z(net_12124) );
SDFF_X2 inst_883 ( .Q(net_8562), .D(net_8562), .SI(net_3947), .SE(net_3878), .CK(net_12407) );
CLKBUF_X2 inst_12536 ( .A(net_12383), .Z(net_12384) );
CLKBUF_X2 inst_12710 ( .A(net_12557), .Z(net_12558) );
SDFF_X2 inst_756 ( .Q(net_8797), .D(net_8797), .SI(net_3974), .SE(net_3879), .CK(net_9993) );
CLKBUF_X2 inst_13423 ( .A(net_13270), .Z(net_13271) );
CLKBUF_X2 inst_9270 ( .A(net_9117), .Z(net_9118) );
CLKBUF_X2 inst_15628 ( .A(net_13007), .Z(net_15476) );
DFFR_X2 inst_7150 ( .QN(net_6486), .D(net_2896), .CK(net_11732), .RN(x6501) );
CLKBUF_X2 inst_15500 ( .A(net_11484), .Z(net_15348) );
CLKBUF_X2 inst_9873 ( .A(net_9373), .Z(net_9721) );
CLKBUF_X2 inst_9685 ( .A(net_9219), .Z(net_9533) );
SDFF_X2 inst_1165 ( .SI(net_7320), .Q(net_6595), .D(net_6595), .SE(net_3069), .CK(net_9835) );
INV_X4 inst_5439 ( .ZN(net_1363), .A(net_822) );
CLKBUF_X2 inst_11029 ( .A(net_9147), .Z(net_10877) );
AOI21_X2 inst_8891 ( .B2(net_5871), .ZN(net_5797), .A(net_5790), .B1(net_2682) );
SDFFR_X1 inst_2644 ( .D(net_6767), .SE(net_4506), .CK(net_9252), .RN(x6501), .SI(x1855), .Q(x1855) );
DFFS_X1 inst_6922 ( .D(net_6145), .CK(net_13660), .SN(x6501), .Q(x794) );
SDFFR_X2 inst_2626 ( .Q(net_7377), .D(net_7377), .SE(net_1136), .CK(net_18620), .RN(x6501), .SI(x4764) );
CLKBUF_X2 inst_9314 ( .A(net_9142), .Z(net_9162) );
NAND2_X2 inst_4629 ( .ZN(net_5452), .A1(net_2946), .A2(net_2518) );
CLKBUF_X2 inst_17307 ( .A(net_17154), .Z(net_17155) );
CLKBUF_X2 inst_14140 ( .A(net_13987), .Z(net_13988) );
INV_X4 inst_5983 ( .A(net_6317), .ZN(net_1254) );
AND2_X4 inst_9056 ( .A1(net_3948), .ZN(net_3901), .A2(net_3277) );
CLKBUF_X2 inst_17629 ( .A(net_17476), .Z(net_17477) );
CLKBUF_X2 inst_16825 ( .A(net_16066), .Z(net_16673) );
DFFS_X2 inst_6883 ( .QN(net_6149), .D(net_3118), .CK(net_18475), .SN(x6501) );
CLKBUF_X2 inst_17107 ( .A(net_16954), .Z(net_16955) );
SDFF_X2 inst_992 ( .D(net_7312), .SI(net_6620), .Q(net_6620), .SE(net_3123), .CK(net_12038) );
CLKBUF_X2 inst_18040 ( .A(net_16053), .Z(net_17888) );
SDFF_X2 inst_488 ( .SI(net_8612), .Q(net_8612), .SE(net_3984), .D(net_3974), .CK(net_10844) );
CLKBUF_X2 inst_14085 ( .A(net_13374), .Z(net_13933) );
AOI22_X2 inst_7809 ( .A2(net_8236), .B2(net_6144), .A1(net_4764), .ZN(net_4756), .B1(net_4522) );
INV_X4 inst_5196 ( .A(net_2963), .ZN(net_2852) );
CLKBUF_X2 inst_18269 ( .A(net_11125), .Z(net_18117) );
AOI222_X1 inst_8666 ( .A2(net_3599), .B2(net_3598), .C2(net_3597), .ZN(net_3592), .C1(net_1645), .A1(net_1357), .B1(net_917) );
DFFR_X2 inst_7308 ( .D(net_7170), .QN(net_7168), .CK(net_9560), .RN(x6501) );
XNOR2_X2 inst_254 ( .A(net_2750), .B(net_2686), .ZN(net_1195) );
INV_X4 inst_6053 ( .A(net_6403), .ZN(net_890) );
CLKBUF_X2 inst_9543 ( .A(net_9087), .Z(net_9391) );
SDFF_X2 inst_1412 ( .Q(net_7116), .D(net_7116), .SE(net_6278), .SI(net_2544), .CK(net_15908) );
CLKBUF_X2 inst_9862 ( .A(net_9709), .Z(net_9710) );
CLKBUF_X2 inst_17066 ( .A(net_16913), .Z(net_16914) );
CLKBUF_X2 inst_10957 ( .A(net_10804), .Z(net_10805) );
CLKBUF_X2 inst_15382 ( .A(net_15229), .Z(net_15230) );
CLKBUF_X2 inst_13364 ( .A(net_13211), .Z(net_13212) );
CLKBUF_X2 inst_12774 ( .A(net_12621), .Z(net_12622) );
SDFF_X2 inst_661 ( .Q(net_8435), .D(net_8435), .SI(net_3941), .SE(net_3934), .CK(net_10354) );
INV_X2 inst_6265 ( .A(net_8245), .ZN(net_4632) );
DFFR_X1 inst_7416 ( .D(net_5673), .CK(net_13900), .RN(x6501), .Q(x563) );
CLKBUF_X2 inst_10817 ( .A(net_10664), .Z(net_10665) );
SDFFS_X2 inst_2073 ( .SI(net_7374), .SE(net_2794), .Q(net_163), .D(net_163), .CK(net_17739), .SN(x6501) );
DFFR_X2 inst_7346 ( .Q(net_7333), .CK(net_11659), .D(x12980), .RN(x6501) );
AOI222_X1 inst_8661 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3905), .B1(net_3275), .C1(net_3274), .A1(x13712) );
CLKBUF_X2 inst_11418 ( .A(net_11265), .Z(net_11266) );
NAND3_X2 inst_3984 ( .A3(net_1894), .ZN(net_1834), .A1(net_1626), .A2(net_272) );
NAND2_X2 inst_4682 ( .A2(net_2161), .ZN(net_2152), .A1(net_2068) );
CLKBUF_X2 inst_17161 ( .A(net_9584), .Z(net_17009) );
CLKBUF_X2 inst_11310 ( .A(net_10101), .Z(net_11158) );
SDFF_X2 inst_419 ( .SI(net_8300), .Q(net_8300), .SE(net_3978), .D(net_3977), .CK(net_11115) );
DFFR_X1 inst_7488 ( .Q(net_8890), .D(net_3904), .CK(net_11270), .RN(x6501) );
CLKBUF_X2 inst_12546 ( .A(net_11535), .Z(net_12394) );
CLKBUF_X2 inst_12098 ( .A(net_11945), .Z(net_11946) );
INV_X2 inst_6495 ( .A(net_8267), .ZN(net_550) );
CLKBUF_X2 inst_15763 ( .A(net_15610), .Z(net_15611) );
DFFS_X1 inst_6941 ( .D(net_6145), .CK(net_13645), .SN(x6501), .Q(x749) );
CLKBUF_X2 inst_18201 ( .A(net_11849), .Z(net_18049) );
CLKBUF_X2 inst_10629 ( .A(net_10476), .Z(net_10477) );
CLKBUF_X2 inst_14298 ( .A(net_14145), .Z(net_14146) );
CLKBUF_X2 inst_14283 ( .A(net_14130), .Z(net_14131) );
CLKBUF_X2 inst_16222 ( .A(net_12114), .Z(net_16070) );
CLKBUF_X2 inst_12377 ( .A(net_10125), .Z(net_12225) );
AOI22_X2 inst_7898 ( .B1(net_8981), .A2(net_5538), .B2(net_5456), .ZN(net_4531), .A1(net_410) );
CLKBUF_X2 inst_16848 ( .A(net_16695), .Z(net_16696) );
CLKBUF_X2 inst_12749 ( .A(net_12596), .Z(net_12597) );
CLKBUF_X2 inst_11160 ( .A(net_11007), .Z(net_11008) );
XOR2_X2 inst_34 ( .B(net_2725), .A(net_2676), .Z(net_1191) );
NAND4_X2 inst_3717 ( .A4(net_6236), .A1(net_6235), .ZN(net_4420), .A2(net_3655), .A3(net_3654) );
AND2_X4 inst_9120 ( .A2(net_9054), .A1(net_2520), .ZN(net_1496) );
XOR2_X2 inst_12 ( .Z(net_1512), .B(net_1511), .A(net_1166) );
CLKBUF_X2 inst_12690 ( .A(net_10733), .Z(net_12538) );
CLKBUF_X2 inst_9823 ( .A(net_9670), .Z(net_9671) );
CLKBUF_X2 inst_13946 ( .A(net_13793), .Z(net_13794) );
CLKBUF_X2 inst_18520 ( .A(net_18367), .Z(net_18368) );
CLKBUF_X2 inst_18674 ( .A(net_18521), .Z(net_18522) );
CLKBUF_X2 inst_9856 ( .A(net_9703), .Z(net_9704) );
SDFF_X2 inst_1424 ( .SI(net_7281), .Q(net_7058), .D(net_7058), .SE(net_6280), .CK(net_19041) );
SDFF_X2 inst_1425 ( .SI(net_7264), .Q(net_7041), .D(net_7041), .SE(net_6280), .CK(net_17088) );
SDFFR_X2 inst_2198 ( .SI(net_6485), .Q(net_6482), .D(net_6482), .SE(net_2897), .CK(net_11701), .RN(x6501) );
XNOR2_X2 inst_258 ( .ZN(net_1189), .A(net_1188), .B(net_883) );
SDFFR_X2 inst_2405 ( .SI(net_7368), .SE(net_2740), .D(net_2693), .QN(net_279), .CK(net_16418), .RN(x6501) );
CLKBUF_X2 inst_13126 ( .A(net_12973), .Z(net_12974) );
OAI21_X2 inst_3076 ( .ZN(net_3883), .B2(net_3552), .A(net_3363), .B1(net_1342) );
CLKBUF_X2 inst_10964 ( .A(net_10541), .Z(net_10812) );
SDFF_X2 inst_482 ( .SI(net_8604), .Q(net_8604), .SE(net_3984), .D(net_3962), .CK(net_10182) );
CLKBUF_X2 inst_9804 ( .A(net_9200), .Z(net_9652) );
CLKBUF_X2 inst_19190 ( .A(net_14597), .Z(net_19038) );
NOR2_X2 inst_3534 ( .ZN(net_4274), .A2(net_1584), .A1(net_1369) );
NOR3_X2 inst_3276 ( .ZN(net_2793), .A1(net_2400), .A3(net_2398), .A2(net_2389) );
CLKBUF_X2 inst_10230 ( .A(net_9598), .Z(net_10078) );
NAND3_X2 inst_3996 ( .ZN(net_4412), .A3(net_4322), .A1(net_1521), .A2(net_1309) );
DFFR_X2 inst_7059 ( .Q(net_6796), .D(net_6259), .CK(net_9578), .RN(x6501) );
SDFF_X2 inst_539 ( .Q(net_8680), .D(net_8680), .SI(net_3966), .SE(net_3935), .CK(net_10938) );
CLKBUF_X2 inst_12915 ( .A(net_12762), .Z(net_12763) );
CLKBUF_X2 inst_11066 ( .A(net_10913), .Z(net_10914) );
SDFF_X2 inst_895 ( .SI(net_8739), .Q(net_8739), .SE(net_6195), .D(net_3949), .CK(net_12576) );
CLKBUF_X2 inst_11042 ( .A(net_10889), .Z(net_10890) );
CLKBUF_X2 inst_10054 ( .A(net_9746), .Z(net_9902) );
INV_X2 inst_6583 ( .A(net_8966), .ZN(net_1648) );
CLKBUF_X2 inst_10034 ( .A(net_9172), .Z(net_9882) );
SDFFR_X2 inst_2341 ( .SI(net_7559), .Q(net_7559), .D(net_2760), .SE(net_2347), .CK(net_13694), .RN(x6501) );
INV_X4 inst_5526 ( .ZN(net_867), .A(net_664) );
CLKBUF_X2 inst_10685 ( .A(net_10229), .Z(net_10533) );
CLKBUF_X2 inst_10616 ( .A(net_10164), .Z(net_10464) );
NAND2_X2 inst_4122 ( .ZN(net_5404), .A2(net_5228), .A1(net_5132) );
CLKBUF_X2 inst_12557 ( .A(net_12404), .Z(net_12405) );
CLKBUF_X2 inst_13184 ( .A(net_13031), .Z(net_13032) );
CLKBUF_X2 inst_9901 ( .A(net_9748), .Z(net_9749) );
CLKBUF_X2 inst_16482 ( .A(net_13391), .Z(net_16330) );
CLKBUF_X2 inst_10324 ( .A(net_10171), .Z(net_10172) );
CLKBUF_X2 inst_16340 ( .A(net_14357), .Z(net_16188) );
AND2_X2 inst_9189 ( .ZN(net_1929), .A1(net_1760), .A2(net_1759) );
NAND2_X2 inst_4797 ( .ZN(net_1439), .A1(net_1112), .A2(net_951) );
INV_X4 inst_6082 ( .A(net_7160), .ZN(net_731) );
AOI22_X2 inst_8482 ( .B1(net_6676), .A1(net_6643), .A2(net_6213), .B2(net_6138), .ZN(net_3458) );
SDFF_X2 inst_826 ( .SI(net_8485), .Q(net_8485), .D(net_3977), .SE(net_3884), .CK(net_13089) );
CLKBUF_X2 inst_9343 ( .A(net_9190), .Z(net_9191) );
CLKBUF_X2 inst_16541 ( .A(net_12428), .Z(net_16389) );
NAND3_X2 inst_4002 ( .ZN(net_2652), .A1(net_1324), .A3(net_1323), .A2(net_607) );
CLKBUF_X2 inst_14009 ( .A(net_13856), .Z(net_13857) );
CLKBUF_X2 inst_10362 ( .A(net_10209), .Z(net_10210) );
XNOR2_X2 inst_159 ( .ZN(net_1851), .B(net_1762), .A(net_1761) );
DFFR_X2 inst_7042 ( .QN(net_7496), .D(net_4877), .CK(net_17252), .RN(x6501) );
CLKBUF_X2 inst_13220 ( .A(net_13067), .Z(net_13068) );
CLKBUF_X2 inst_18680 ( .A(net_18527), .Z(net_18528) );
CLKBUF_X2 inst_9572 ( .A(net_9419), .Z(net_9420) );
CLKBUF_X2 inst_15281 ( .A(net_15128), .Z(net_15129) );
INV_X4 inst_5759 ( .A(net_7520), .ZN(net_740) );
CLKBUF_X2 inst_13657 ( .A(net_13504), .Z(net_13505) );
CLKBUF_X2 inst_11005 ( .A(net_9456), .Z(net_10853) );
INV_X2 inst_6318 ( .ZN(net_3345), .A(net_3290) );
DFFR_X1 inst_7379 ( .D(net_5893), .CK(net_11445), .RN(x6501), .Q(x2451) );
CLKBUF_X2 inst_15491 ( .A(net_14414), .Z(net_15339) );
AOI22_X2 inst_8339 ( .A1(net_8625), .B1(net_8440), .A2(net_3864), .B2(net_3863), .ZN(net_3708) );
XOR2_X2 inst_19 ( .Z(net_1414), .B(net_1413), .A(net_921) );
CLKBUF_X2 inst_13623 ( .A(net_12805), .Z(net_13471) );
CLKBUF_X2 inst_11509 ( .A(net_11356), .Z(net_11357) );
CLKBUF_X2 inst_10378 ( .A(net_9811), .Z(net_10226) );
CLKBUF_X2 inst_13599 ( .A(net_13446), .Z(net_13447) );
NAND2_X2 inst_4268 ( .A1(net_7036), .A2(net_5249), .ZN(net_5192) );
CLKBUF_X2 inst_18487 ( .A(net_15652), .Z(net_18335) );
CLKBUF_X2 inst_14170 ( .A(net_9697), .Z(net_14018) );
NAND4_X2 inst_3830 ( .ZN(net_2471), .A4(net_2406), .A1(net_1725), .A3(net_1608), .A2(net_1607) );
CLKBUF_X2 inst_16706 ( .A(net_16553), .Z(net_16554) );
CLKBUF_X2 inst_12287 ( .A(net_12134), .Z(net_12135) );
SDFF_X2 inst_1686 ( .Q(net_8169), .D(net_8169), .SI(net_2749), .SE(net_2538), .CK(net_13755) );
CLKBUF_X2 inst_10541 ( .A(net_9685), .Z(net_10389) );
CLKBUF_X2 inst_15732 ( .A(net_12344), .Z(net_15580) );
CLKBUF_X2 inst_16724 ( .A(net_16571), .Z(net_16572) );
SDFF_X2 inst_1789 ( .D(net_7269), .SI(net_7006), .Q(net_7006), .SE(net_6277), .CK(net_16811) );
CLKBUF_X2 inst_14664 ( .A(net_14314), .Z(net_14512) );
DFFR_X2 inst_7192 ( .QN(net_7225), .D(net_2448), .CK(net_15197), .RN(x6501) );
CLKBUF_X2 inst_14832 ( .A(net_10315), .Z(net_14680) );
CLKBUF_X2 inst_15803 ( .A(net_15650), .Z(net_15651) );
CLKBUF_X2 inst_15951 ( .A(net_11831), .Z(net_15799) );
CLKBUF_X2 inst_18251 ( .A(net_13290), .Z(net_18099) );
CLKBUF_X2 inst_9437 ( .A(net_9284), .Z(net_9285) );
NOR2_X2 inst_3441 ( .A2(net_3093), .ZN(net_3054), .A1(net_2824) );
DFFS_X1 inst_6955 ( .D(net_3231), .CK(net_16331), .SN(x6501), .Q(x905) );
CLKBUF_X2 inst_12332 ( .A(net_12179), .Z(net_12180) );
CLKBUF_X2 inst_9413 ( .A(net_9260), .Z(net_9261) );
AOI22_X2 inst_8000 ( .B1(net_8199), .A1(net_7689), .B2(net_6099), .A2(net_4399), .ZN(net_4133) );
CLKBUF_X2 inst_11535 ( .A(net_11283), .Z(net_11383) );
CLKBUF_X2 inst_15250 ( .A(net_15097), .Z(net_15098) );
CLKBUF_X2 inst_17865 ( .A(net_17712), .Z(net_17713) );
CLKBUF_X2 inst_16715 ( .A(net_16562), .Z(net_16563) );
CLKBUF_X2 inst_12516 ( .A(net_12363), .Z(net_12364) );
CLKBUF_X2 inst_17791 ( .A(net_12672), .Z(net_17639) );
NAND2_X2 inst_4860 ( .ZN(net_2097), .A2(net_567), .A1(net_566) );
CLKBUF_X2 inst_14923 ( .A(net_14593), .Z(net_14771) );
CLKBUF_X2 inst_12226 ( .A(net_9851), .Z(net_12074) );
DFF_X1 inst_6770 ( .Q(net_7549), .D(net_4602), .CK(net_12768) );
CLKBUF_X2 inst_16314 ( .A(net_16161), .Z(net_16162) );
SDFF_X2 inst_1344 ( .Q(net_8195), .D(net_8195), .SI(net_2576), .SE(net_2561), .CK(net_16072) );
SDFF_X2 inst_1460 ( .SI(net_7281), .Q(net_7138), .D(net_7138), .SE(net_6279), .CK(net_19035) );
SDFFR_X2 inst_2287 ( .SI(net_8901), .Q(net_8901), .SE(net_6117), .D(net_2407), .CK(net_16254), .RN(x6501) );
CLKBUF_X2 inst_17336 ( .A(net_14175), .Z(net_17184) );
AOI21_X2 inst_8968 ( .B2(net_6264), .A(net_6151), .ZN(net_2990), .B1(net_1638) );
SDFFR_X2 inst_2630 ( .Q(net_7379), .D(net_7379), .SE(net_1136), .CK(net_18610), .RN(x6501), .SI(x4743) );
CLKBUF_X2 inst_15422 ( .A(net_15269), .Z(net_15270) );
CLKBUF_X2 inst_17329 ( .A(net_17176), .Z(net_17177) );
CLKBUF_X2 inst_17611 ( .A(net_17458), .Z(net_17459) );
SDFF_X2 inst_1443 ( .SI(net_7289), .Q(net_7106), .D(net_7106), .SE(net_6278), .CK(net_18401) );
SDFF_X2 inst_1028 ( .SI(net_7338), .Q(net_6745), .D(net_6745), .SE(net_3124), .CK(net_9486) );
INV_X4 inst_5891 ( .A(net_7613), .ZN(net_807) );
CLKBUF_X2 inst_10107 ( .A(net_9954), .Z(net_9955) );
NAND3_X2 inst_3935 ( .ZN(net_5515), .A1(net_5277), .A2(net_4655), .A3(net_4566) );
CLKBUF_X2 inst_9645 ( .A(net_9462), .Z(net_9493) );
SDFF_X2 inst_1271 ( .Q(net_7811), .D(net_7811), .SE(net_2730), .SI(net_2659), .CK(net_15469) );
CLKBUF_X2 inst_12110 ( .A(net_10576), .Z(net_11958) );
SDFFR_X2 inst_2321 ( .D(net_3388), .SE(net_2685), .SI(net_426), .Q(net_426), .CK(net_17284), .RN(x6501) );
CLKBUF_X2 inst_17503 ( .A(net_17350), .Z(net_17351) );
CLKBUF_X2 inst_13927 ( .A(net_13774), .Z(net_13775) );
CLKBUF_X2 inst_9928 ( .A(net_9775), .Z(net_9776) );
NAND2_X2 inst_4425 ( .A1(net_6863), .A2(net_5016), .ZN(net_5002) );
CLKBUF_X2 inst_9727 ( .A(net_9425), .Z(net_9575) );
NAND2_X2 inst_4461 ( .ZN(net_4907), .A2(net_4694), .A1(net_4533) );
INV_X16 inst_6626 ( .ZN(net_4400), .A(net_3558) );
CLKBUF_X2 inst_14332 ( .A(net_14179), .Z(net_14180) );
DFFR_X1 inst_7407 ( .D(net_5705), .CK(net_17166), .RN(x6501), .Q(x364) );
CLKBUF_X2 inst_12343 ( .A(net_9827), .Z(net_12191) );
CLKBUF_X2 inst_10807 ( .A(net_10654), .Z(net_10655) );
CLKBUF_X2 inst_17221 ( .A(net_17068), .Z(net_17069) );
SDFFR_X2 inst_2236 ( .Q(net_7460), .D(net_7460), .SE(net_2863), .CK(net_10626), .SI(x13508), .RN(x6501) );
NOR2_X2 inst_3368 ( .ZN(net_5557), .A2(net_5356), .A1(net_5355) );
DFFR_X2 inst_7307 ( .QN(net_8270), .D(net_8266), .CK(net_15651), .RN(x6501) );
SDFF_X2 inst_1553 ( .Q(net_7981), .D(net_7981), .SI(net_2659), .SE(net_2542), .CK(net_15527) );
CLKBUF_X2 inst_13038 ( .A(net_12885), .Z(net_12886) );
CLKBUF_X2 inst_13937 ( .A(net_13784), .Z(net_13785) );
CLKBUF_X2 inst_16027 ( .A(net_13130), .Z(net_15875) );
CLKBUF_X2 inst_15322 ( .A(net_13986), .Z(net_15170) );
CLKBUF_X2 inst_10458 ( .A(net_10305), .Z(net_10306) );
SDFF_X2 inst_1635 ( .Q(net_8150), .D(net_8150), .SI(net_2709), .SE(net_2538), .CK(net_15759) );
NAND2_X2 inst_4130 ( .ZN(net_5393), .A1(net_5223), .A2(net_5004) );
CLKBUF_X2 inst_12121 ( .A(net_11968), .Z(net_11969) );
CLKBUF_X2 inst_13102 ( .A(net_12949), .Z(net_12950) );
CLKBUF_X2 inst_17515 ( .A(net_13180), .Z(net_17363) );
SDFF_X2 inst_1500 ( .SI(net_7858), .Q(net_7858), .D(net_2590), .SE(net_2558), .CK(net_15999) );
CLKBUF_X2 inst_14737 ( .A(net_14584), .Z(net_14585) );
CLKBUF_X2 inst_11731 ( .A(net_11578), .Z(net_11579) );
OR3_X2 inst_2805 ( .ZN(net_4410), .A3(net_4406), .A1(net_4390), .A2(net_4380) );
INV_X2 inst_6438 ( .ZN(net_816), .A(net_642) );
OAI22_X2 inst_2932 ( .B2(net_2299), .A2(net_2187), .ZN(net_2178), .A1(net_2177), .B1(net_1472) );
CLKBUF_X2 inst_17891 ( .A(net_17738), .Z(net_17739) );
CLKBUF_X2 inst_18329 ( .A(net_13413), .Z(net_18177) );
DFFS_X1 inst_6917 ( .Q(net_7162), .D(net_4625), .CK(net_9549), .SN(x6501) );
CLKBUF_X2 inst_17581 ( .A(net_17428), .Z(net_17429) );
CLKBUF_X2 inst_9483 ( .A(net_9330), .Z(net_9331) );
CLKBUF_X2 inst_15839 ( .A(net_15686), .Z(net_15687) );
OAI21_X2 inst_3048 ( .B2(net_8229), .B1(net_4850), .ZN(net_4763), .A(net_2617) );
CLKBUF_X2 inst_10911 ( .A(net_10758), .Z(net_10759) );
NAND2_X2 inst_4854 ( .A2(net_8893), .A1(net_3000), .ZN(net_1423) );
CLKBUF_X2 inst_13862 ( .A(net_13709), .Z(net_13710) );
NOR2_X2 inst_3346 ( .ZN(net_5579), .A1(net_5446), .A2(net_5445) );
OAI21_X2 inst_2992 ( .B2(net_5912), .ZN(net_5901), .A(net_5800), .B1(net_1124) );
SDFF_X2 inst_1080 ( .D(net_7331), .SI(net_6507), .Q(net_6507), .SE(net_3071), .CK(net_9064) );
INV_X2 inst_6405 ( .A(net_6418), .ZN(net_1079) );
SDFFR_X2 inst_2374 ( .SE(net_2260), .Q(net_320), .D(net_320), .CK(net_10434), .RN(x6501), .SI(x3122) );
DFFR_X1 inst_7473 ( .QN(net_7424), .D(net_4215), .CK(net_12393), .RN(x6501) );
CLKBUF_X2 inst_15723 ( .A(net_15570), .Z(net_15571) );
SDFF_X2 inst_1103 ( .D(net_7333), .SI(net_6542), .Q(net_6542), .SE(net_3086), .CK(net_11674) );
INV_X2 inst_6535 ( .A(net_8951), .ZN(net_519) );
AOI222_X1 inst_8620 ( .A2(net_8224), .A1(net_4891), .B2(net_4889), .C2(net_4888), .ZN(net_4886), .C1(net_3131), .B1(net_2669) );
CLKBUF_X2 inst_17709 ( .A(net_17556), .Z(net_17557) );
CLKBUF_X2 inst_10678 ( .A(net_10347), .Z(net_10526) );
CLKBUF_X2 inst_9256 ( .A(net_9074), .Z(net_9104) );
DFFR_X1 inst_7494 ( .D(net_3209), .CK(net_16522), .RN(x6501), .Q(x43) );
SDFF_X2 inst_549 ( .Q(net_8694), .D(net_8694), .SI(net_3941), .SE(net_3935), .CK(net_12895) );
NAND2_X2 inst_4329 ( .A1(net_7141), .A2(net_5166), .ZN(net_5128) );
CLKBUF_X2 inst_12566 ( .A(net_12413), .Z(net_12414) );
NAND2_X2 inst_4708 ( .ZN(net_2659), .A2(net_1586), .A1(net_1121) );
CLKBUF_X2 inst_18886 ( .A(net_18733), .Z(net_18734) );
INV_X4 inst_5202 ( .ZN(net_5843), .A(net_5718) );
CLKBUF_X2 inst_13617 ( .A(net_13464), .Z(net_13465) );
INV_X2 inst_6231 ( .ZN(net_5479), .A(net_5302) );
CLKBUF_X2 inst_19084 ( .A(net_18931), .Z(net_18932) );
CLKBUF_X2 inst_16592 ( .A(net_11000), .Z(net_16440) );
CLKBUF_X2 inst_16539 ( .A(net_16386), .Z(net_16387) );
CLKBUF_X2 inst_13776 ( .A(net_13623), .Z(net_13624) );
INV_X2 inst_6331 ( .A(net_5830), .ZN(net_3060) );
CLKBUF_X2 inst_16962 ( .A(net_16809), .Z(net_16810) );
CLKBUF_X2 inst_9737 ( .A(net_9584), .Z(net_9585) );
SDFFR_X1 inst_2673 ( .SI(net_7527), .SE(net_5043), .CK(net_11951), .RN(x6501), .Q(x4214), .D(x4214) );
CLKBUF_X2 inst_13592 ( .A(net_13439), .Z(net_13440) );
SDFF_X2 inst_1618 ( .Q(net_8160), .D(net_8160), .SI(net_2589), .SE(net_2538), .CK(net_18369) );
INV_X4 inst_5062 ( .ZN(net_5938), .A(net_5936) );
CLKBUF_X2 inst_14166 ( .A(net_14013), .Z(net_14014) );
SDFFR_X2 inst_2126 ( .SI(net_7191), .Q(net_7191), .D(net_6442), .SE(net_4362), .CK(net_16264), .RN(x6501) );
CLKBUF_X2 inst_10484 ( .A(net_10331), .Z(net_10332) );
CLKBUF_X2 inst_18917 ( .A(net_18764), .Z(net_18765) );
AOI22_X2 inst_7776 ( .B1(net_6966), .A1(net_6926), .A2(net_5443), .B2(net_5442), .ZN(net_5299) );
SDFFR_X1 inst_2765 ( .QN(net_7582), .D(net_3956), .SE(net_3144), .SI(net_749), .CK(net_11035), .RN(x6501) );
NOR2_X2 inst_3600 ( .A1(net_1076), .ZN(net_842), .A2(net_546) );
XNOR2_X2 inst_219 ( .ZN(net_1404), .B(net_1403), .A(net_712) );
NAND2_X2 inst_4881 ( .A2(net_7392), .ZN(net_776), .A1(net_181) );
CLKBUF_X2 inst_15320 ( .A(net_15167), .Z(net_15168) );
AOI21_X2 inst_8980 ( .B2(net_2077), .ZN(net_2059), .A(net_1927), .B1(net_1777) );
INV_X4 inst_5501 ( .ZN(net_1633), .A(net_701) );
SDFFR_X2 inst_2204 ( .SI(net_9052), .Q(net_9052), .SE(net_2963), .D(net_2235), .CK(net_11196), .RN(x6501) );
CLKBUF_X2 inst_16785 ( .A(net_15052), .Z(net_16633) );
CLKBUF_X2 inst_16595 ( .A(net_12353), .Z(net_16443) );
SDFF_X2 inst_1609 ( .Q(net_8115), .D(net_8115), .SI(net_2655), .SE(net_2541), .CK(net_15435) );
NAND2_X2 inst_4105 ( .ZN(net_5427), .A2(net_5240), .A1(net_5150) );
CLKBUF_X2 inst_16530 ( .A(net_16377), .Z(net_16378) );
CLKBUF_X2 inst_16984 ( .A(net_13926), .Z(net_16832) );
SDFF_X2 inst_408 ( .SI(net_8322), .Q(net_8322), .SE(net_3978), .D(net_3954), .CK(net_10085) );
NAND2_X2 inst_4701 ( .ZN(net_2180), .A2(net_2046), .A1(net_1614) );
INV_X4 inst_5644 ( .A(net_7570), .ZN(net_2969) );
CLKBUF_X2 inst_12419 ( .A(net_12266), .Z(net_12267) );
CLKBUF_X2 inst_11212 ( .A(net_11059), .Z(net_11060) );
CLKBUF_X2 inst_16524 ( .A(net_16371), .Z(net_16372) );
INV_X4 inst_5596 ( .A(net_7584), .ZN(net_594) );
CLKBUF_X2 inst_17374 ( .A(net_17221), .Z(net_17222) );
CLKBUF_X2 inst_11591 ( .A(net_11438), .Z(net_11439) );
CLKBUF_X2 inst_10719 ( .A(net_10478), .Z(net_10567) );
NAND4_X2 inst_3814 ( .ZN(net_3612), .A1(net_3431), .A2(net_3430), .A3(net_3429), .A4(net_3428) );
CLKBUF_X2 inst_12968 ( .A(net_12815), .Z(net_12816) );
AOI22_X2 inst_8498 ( .B1(net_6680), .A1(net_6647), .A2(net_6213), .B2(net_6138), .ZN(net_3442) );
CLKBUF_X2 inst_15605 ( .A(net_15452), .Z(net_15453) );
AOI22_X2 inst_7871 ( .A2(net_6436), .A1(net_5654), .B2(net_4881), .ZN(net_4570), .B1(net_236) );
NOR2_X2 inst_3514 ( .ZN(net_2344), .A1(net_2318), .A2(net_1773) );
CLKBUF_X2 inst_10826 ( .A(net_10302), .Z(net_10674) );
SDFF_X2 inst_1510 ( .SI(net_7871), .Q(net_7871), .D(net_2716), .SE(net_2558), .CK(net_14281) );
XNOR2_X2 inst_121 ( .ZN(net_2983), .A(net_2830), .B(net_1053) );
CLKBUF_X2 inst_16659 ( .A(net_16506), .Z(net_16507) );
CLKBUF_X2 inst_12449 ( .A(net_12296), .Z(net_12297) );
SDFF_X2 inst_1065 ( .D(net_7327), .SI(net_6536), .Q(net_6536), .SE(net_3086), .CK(net_9857) );
CLKBUF_X2 inst_12002 ( .A(net_11849), .Z(net_11850) );
NAND2_X2 inst_4119 ( .ZN(net_5408), .A1(net_5137), .A2(net_5136) );
NAND2_X2 inst_4332 ( .A1(net_7142), .A2(net_5166), .ZN(net_5125) );
CLKBUF_X2 inst_13766 ( .A(net_13613), .Z(net_13614) );
CLKBUF_X2 inst_14348 ( .A(net_11681), .Z(net_14196) );
CLKBUF_X2 inst_9495 ( .A(net_9065), .Z(net_9343) );
INV_X4 inst_5353 ( .A(net_1922), .ZN(net_1176) );
CLKBUF_X2 inst_14189 ( .A(net_14036), .Z(net_14037) );
CLKBUF_X2 inst_9981 ( .A(net_9828), .Z(net_9829) );
CLKBUF_X2 inst_16981 ( .A(net_11096), .Z(net_16829) );
NAND2_X2 inst_4671 ( .ZN(net_2196), .A1(net_2133), .A2(net_1926) );
CLKBUF_X2 inst_16860 ( .A(net_16707), .Z(net_16708) );
SDFF_X2 inst_530 ( .Q(net_8887), .D(net_8887), .SI(net_3949), .SE(net_3936), .CK(net_10571) );
AOI211_X2 inst_9009 ( .C2(net_6431), .C1(net_5654), .ZN(net_5451), .B(net_4955), .A(net_4907) );
AOI22_X2 inst_8004 ( .B1(net_8113), .A1(net_7875), .A2(net_6098), .B2(net_4190), .ZN(net_4130) );
CLKBUF_X2 inst_18417 ( .A(net_10555), .Z(net_18265) );
CLKBUF_X2 inst_18994 ( .A(net_11394), .Z(net_18842) );
SDFF_X2 inst_1353 ( .Q(net_8206), .D(net_8206), .SI(net_2710), .SE(net_2561), .CK(net_13787) );
DFFR_X1 inst_7370 ( .D(net_5930), .CK(net_13910), .RN(x6501), .Q(x626) );
CLKBUF_X2 inst_15483 ( .A(net_15330), .Z(net_15331) );
SDFF_X2 inst_769 ( .Q(net_8813), .D(net_8813), .SI(net_3949), .SE(net_3879), .CK(net_10521) );
CLKBUF_X2 inst_13334 ( .A(net_13181), .Z(net_13182) );
CLKBUF_X2 inst_12429 ( .A(net_12276), .Z(net_12277) );
SDFF_X2 inst_1200 ( .D(net_7300), .SI(net_7037), .Q(net_7037), .SE(net_6277), .CK(net_18220) );
CLKBUF_X2 inst_15593 ( .A(net_15440), .Z(net_15441) );
CLKBUF_X2 inst_10888 ( .A(net_10735), .Z(net_10736) );
CLKBUF_X2 inst_10120 ( .A(net_9967), .Z(net_9968) );
CLKBUF_X2 inst_17001 ( .A(net_16689), .Z(net_16849) );
CLKBUF_X2 inst_15473 ( .A(net_15320), .Z(net_15321) );
CLKBUF_X2 inst_10918 ( .A(net_10765), .Z(net_10766) );
AOI22_X2 inst_8523 ( .B1(net_6589), .A1(net_6556), .A2(net_6257), .B2(net_6110), .ZN(net_3417) );
OAI21_X2 inst_3021 ( .B2(net_5044), .ZN(net_5039), .A(net_4883), .B1(net_2142) );
INV_X2 inst_6349 ( .ZN(net_2350), .A(net_2349) );
CLKBUF_X2 inst_16037 ( .A(net_15884), .Z(net_15885) );
DFFR_X2 inst_7365 ( .Q(net_7321), .CK(net_11358), .D(x13086), .RN(x6501) );
INV_X2 inst_6474 ( .ZN(net_849), .A(net_226) );
CLKBUF_X2 inst_12232 ( .A(net_12079), .Z(net_12080) );
CLKBUF_X2 inst_11664 ( .A(net_11511), .Z(net_11512) );
CLKBUF_X2 inst_15084 ( .A(net_14931), .Z(net_14932) );
CLKBUF_X2 inst_18794 ( .A(net_18641), .Z(net_18642) );
CLKBUF_X2 inst_12618 ( .A(net_12465), .Z(net_12466) );
CLKBUF_X2 inst_13045 ( .A(net_12892), .Z(net_12893) );
CLKBUF_X2 inst_18628 ( .A(net_9612), .Z(net_18476) );
CLKBUF_X2 inst_11922 ( .A(net_11769), .Z(net_11770) );
CLKBUF_X2 inst_14790 ( .A(net_11973), .Z(net_14638) );
NAND3_X2 inst_3911 ( .ZN(net_5627), .A1(net_5556), .A3(net_5490), .A2(net_5350) );
SDFF_X2 inst_1515 ( .SI(net_7849), .Q(net_7849), .D(net_2573), .SE(net_2558), .CK(net_18056) );
DFF_X1 inst_6777 ( .Q(net_7556), .D(net_4595), .CK(net_10474) );
CLKBUF_X2 inst_9743 ( .A(net_9264), .Z(net_9591) );
DFFR_X1 inst_7546 ( .Q(net_6479), .D(net_980), .CK(net_11733), .RN(x6501) );
CLKBUF_X2 inst_13088 ( .A(net_12576), .Z(net_12936) );
SDFF_X2 inst_1782 ( .D(net_7265), .SI(net_6962), .Q(net_6962), .SE(net_6283), .CK(net_17425) );
CLKBUF_X2 inst_15274 ( .A(net_15121), .Z(net_15122) );
NAND2_X2 inst_4472 ( .A2(net_5463), .ZN(net_4645), .A1(net_439) );
DFFR_X1 inst_7513 ( .D(net_6417), .Q(net_6408), .CK(net_9677), .RN(x6501) );
SDFF_X2 inst_1015 ( .SI(net_7330), .Q(net_6671), .D(net_6671), .SE(net_3126), .CK(net_11331) );
CLKBUF_X2 inst_15776 ( .A(net_15623), .Z(net_15624) );
DFFR_X2 inst_7003 ( .D(net_5881), .CK(net_11485), .RN(x6501), .Q(x2400) );
CLKBUF_X2 inst_14390 ( .A(net_12437), .Z(net_14238) );
NAND3_X2 inst_3899 ( .ZN(net_5639), .A1(net_5568), .A3(net_5502), .A2(net_5398) );
CLKBUF_X2 inst_15940 ( .A(net_11368), .Z(net_15788) );
CLKBUF_X2 inst_14226 ( .A(net_14073), .Z(net_14074) );
OAI211_X2 inst_3213 ( .B(net_2304), .ZN(net_1909), .C2(net_1908), .A(net_1292), .C1(net_666) );
CLKBUF_X2 inst_17254 ( .A(net_11529), .Z(net_17102) );
CLKBUF_X2 inst_15771 ( .A(net_15618), .Z(net_15619) );
SDFF_X2 inst_1661 ( .SI(net_7753), .Q(net_7753), .D(net_2576), .SE(net_2560), .CK(net_16035) );
CLKBUF_X2 inst_13583 ( .A(net_12474), .Z(net_13431) );
XNOR2_X2 inst_283 ( .A(net_2137), .B(net_1778), .ZN(net_1015) );
CLKBUF_X2 inst_15193 ( .A(net_15040), .Z(net_15041) );
SDFFR_X2 inst_2519 ( .Q(net_6421), .D(net_6421), .SE(net_2433), .SI(net_1146), .CK(net_18658), .RN(x6501) );
NOR2_X2 inst_3406 ( .ZN(net_4554), .A2(net_3578), .A1(net_1708) );
SDFF_X2 inst_1597 ( .Q(net_8113), .D(net_8113), .SI(net_2585), .SE(net_2541), .CK(net_15826) );
DFFR_X1 inst_7574 ( .Q(net_8286), .D(net_8276), .CK(net_12227), .RN(x6501) );
CLKBUF_X2 inst_18000 ( .A(net_17847), .Z(net_17848) );
CLKBUF_X2 inst_18951 ( .A(net_16015), .Z(net_18799) );
SDFF_X2 inst_431 ( .Q(net_8759), .D(net_8759), .SE(net_3982), .SI(net_3958), .CK(net_10028) );
INV_X4 inst_6063 ( .A(net_7505), .ZN(net_4457) );
CLKBUF_X2 inst_11331 ( .A(net_11178), .Z(net_11179) );
DFFS_X2 inst_6906 ( .QN(net_8267), .D(net_8263), .CK(net_18466), .SN(x6501) );
DFFR_X1 inst_7429 ( .QN(net_8930), .D(net_4858), .CK(net_17326), .RN(x6501) );
CLKBUF_X2 inst_15657 ( .A(net_11285), .Z(net_15505) );
SDFF_X2 inst_1364 ( .Q(net_8184), .D(net_8184), .SI(net_2709), .SE(net_2561), .CK(net_18557) );
CLKBUF_X2 inst_11514 ( .A(net_11361), .Z(net_11362) );
CLKBUF_X2 inst_18105 ( .A(net_13290), .Z(net_17953) );
CLKBUF_X2 inst_14460 ( .A(net_14307), .Z(net_14308) );
DFF_X1 inst_6847 ( .Q(net_6435), .D(net_3634), .CK(net_17958) );
CLKBUF_X2 inst_16417 ( .A(net_15282), .Z(net_16265) );
CLKBUF_X2 inst_14563 ( .A(net_14410), .Z(net_14411) );
CLKBUF_X2 inst_14801 ( .A(net_14648), .Z(net_14649) );
CLKBUF_X2 inst_11278 ( .A(net_11125), .Z(net_11126) );
CLKBUF_X2 inst_18366 ( .A(net_18213), .Z(net_18214) );
CLKBUF_X2 inst_9560 ( .A(net_9196), .Z(net_9408) );
SDFFR_X2 inst_2544 ( .QN(net_6366), .SE(net_2147), .SI(net_1942), .D(net_966), .CK(net_14753), .RN(x6501) );
CLKBUF_X2 inst_15329 ( .A(net_15176), .Z(net_15177) );
CLKBUF_X2 inst_19118 ( .A(net_17156), .Z(net_18966) );
CLKBUF_X2 inst_16854 ( .A(net_16701), .Z(net_16702) );
CLKBUF_X2 inst_14364 ( .A(net_11740), .Z(net_14212) );
SDFF_X2 inst_685 ( .Q(net_8683), .D(net_8683), .SI(net_3944), .SE(net_3935), .CK(net_12265) );
CLKBUF_X2 inst_13281 ( .A(net_13128), .Z(net_13129) );
CLKBUF_X2 inst_9586 ( .A(net_9433), .Z(net_9434) );
CLKBUF_X2 inst_15478 ( .A(net_15325), .Z(net_15326) );
CLKBUF_X2 inst_15236 ( .A(net_15083), .Z(net_15084) );
CLKBUF_X2 inst_13829 ( .A(net_13676), .Z(net_13677) );
CLKBUF_X2 inst_17485 ( .A(net_15453), .Z(net_17333) );
AND2_X4 inst_9150 ( .ZN(net_6279), .A2(net_2265), .A1(net_1427) );
INV_X2 inst_6338 ( .ZN(net_2856), .A(net_2788) );
INV_X2 inst_6561 ( .A(net_8967), .ZN(net_1927) );
CLKBUF_X2 inst_12700 ( .A(net_12547), .Z(net_12548) );
CLKBUF_X2 inst_12678 ( .A(net_12525), .Z(net_12526) );
DFFS_X2 inst_6886 ( .QN(net_8892), .D(net_3001), .CK(net_18923), .SN(x6501) );
SDFF_X2 inst_427 ( .Q(net_8754), .D(net_8754), .SE(net_3982), .SI(net_3966), .CK(net_10033) );
CLKBUF_X2 inst_18592 ( .A(net_18439), .Z(net_18440) );
CLKBUF_X2 inst_13113 ( .A(net_12960), .Z(net_12961) );
CLKBUF_X2 inst_11952 ( .A(net_10668), .Z(net_11800) );
SDFFR_X2 inst_2144 ( .SI(net_7183), .Q(net_7183), .D(net_6434), .SE(net_4362), .CK(net_13725), .RN(x6501) );
CLKBUF_X2 inst_15327 ( .A(net_11642), .Z(net_15175) );
INV_X4 inst_5721 ( .A(net_7251), .ZN(net_1954) );
INV_X4 inst_6121 ( .A(net_5971), .ZN(x3327) );
XNOR2_X2 inst_138 ( .B(net_6321), .ZN(net_2536), .A(net_2535) );
DFF_X1 inst_6793 ( .QN(net_8240), .D(net_4440), .CK(net_14463) );
OR3_X2 inst_2810 ( .A2(net_9004), .ZN(net_1924), .A3(net_1923), .A1(net_1868) );
CLKBUF_X2 inst_16969 ( .A(net_10810), .Z(net_16817) );
SDFF_X2 inst_899 ( .SI(net_8715), .Q(net_8715), .SE(net_6195), .D(net_3962), .CK(net_10126) );
CLKBUF_X2 inst_12304 ( .A(net_12151), .Z(net_12152) );
CLKBUF_X2 inst_13346 ( .A(net_13193), .Z(net_13194) );
CLKBUF_X2 inst_13256 ( .A(net_10697), .Z(net_13104) );
CLKBUF_X2 inst_9889 ( .A(net_9736), .Z(net_9737) );
SDFFR_X2 inst_2149 ( .Q(net_8272), .D(net_8272), .SI(net_6153), .SE(net_2996), .CK(net_18457), .RN(x6501) );
AOI22_X2 inst_8356 ( .A1(net_8628), .B1(net_8443), .A2(net_3864), .B2(net_3863), .ZN(net_3692) );
DFFR_X2 inst_6980 ( .D(net_5906), .CK(net_9343), .RN(x6501), .Q(x3651) );
MUX2_X2 inst_5001 ( .S(net_8901), .A(net_8251), .Z(net_2787), .B(net_1173) );
CLKBUF_X2 inst_11875 ( .A(net_9515), .Z(net_11723) );
CLKBUF_X2 inst_17003 ( .A(net_16850), .Z(net_16851) );
CLKBUF_X2 inst_14470 ( .A(net_14317), .Z(net_14318) );
DFFR_X1 inst_7386 ( .D(net_5848), .CK(net_16784), .RN(x6501), .Q(x451) );
CLKBUF_X2 inst_9950 ( .A(net_9614), .Z(net_9798) );
CLKBUF_X2 inst_9319 ( .A(net_9166), .Z(net_9167) );
AOI22_X2 inst_8172 ( .B1(net_8677), .A1(net_8640), .B2(net_6109), .ZN(net_3858), .A2(net_3857) );
CLKBUF_X2 inst_13899 ( .A(net_13746), .Z(net_13747) );
AOI21_X2 inst_8876 ( .B2(net_5871), .ZN(net_5869), .A(net_5865), .B1(net_2758) );
NAND2_X2 inst_4078 ( .A2(net_6780), .A1(net_5835), .ZN(net_5768) );
NAND2_X2 inst_4067 ( .A2(net_6342), .ZN(net_5884), .A1(net_5738) );
CLKBUF_X2 inst_18846 ( .A(net_15418), .Z(net_18694) );
AND2_X4 inst_9109 ( .ZN(net_2082), .A2(net_1881), .A1(net_1309) );
AOI21_X2 inst_8894 ( .B2(net_5871), .ZN(net_5792), .A(net_5785), .B1(x608) );
CLKBUF_X2 inst_10175 ( .A(net_9670), .Z(net_10023) );
CLKBUF_X2 inst_14972 ( .A(net_14819), .Z(net_14820) );
CLKBUF_X2 inst_14180 ( .A(net_11328), .Z(net_14028) );
AOI21_X2 inst_8885 ( .B2(net_5871), .ZN(net_5813), .A(net_5809), .B1(x434) );
NAND3_X2 inst_3883 ( .ZN(net_5888), .A3(net_5776), .A1(net_4963), .A2(net_4784) );
CLKBUF_X2 inst_10020 ( .A(net_9867), .Z(net_9868) );
CLKBUF_X2 inst_11811 ( .A(net_11658), .Z(net_11659) );
CLKBUF_X2 inst_13451 ( .A(net_12122), .Z(net_13299) );
AND2_X4 inst_9096 ( .ZN(net_2541), .A1(net_2274), .A2(net_2267) );
INV_X4 inst_5818 ( .A(net_8965), .ZN(net_1887) );
INV_X4 inst_5510 ( .A(net_1258), .ZN(net_688) );
DFFR_X2 inst_7041 ( .QN(net_7509), .D(net_4912), .CK(net_14502), .RN(x6501) );
AOI22_X2 inst_8415 ( .B1(net_8676), .A1(net_8639), .B2(net_6109), .A2(net_3857), .ZN(net_3637) );
CLKBUF_X2 inst_12632 ( .A(net_12479), .Z(net_12480) );
CLKBUF_X2 inst_10308 ( .A(net_10155), .Z(net_10156) );
SDFFR_X2 inst_2577 ( .D(net_7389), .QN(net_7249), .SI(net_1959), .SE(net_1379), .CK(net_18120), .RN(x6501) );
CLKBUF_X2 inst_15319 ( .A(net_15166), .Z(net_15167) );
DFFR_X1 inst_7565 ( .D(net_6830), .Q(net_6803), .CK(net_9661), .RN(x6501) );
CLKBUF_X2 inst_16571 ( .A(net_11067), .Z(net_16419) );
CLKBUF_X2 inst_17886 ( .A(net_14947), .Z(net_17734) );
CLKBUF_X2 inst_13267 ( .A(net_13114), .Z(net_13115) );
INV_X2 inst_6431 ( .ZN(net_698), .A(net_697) );
CLKBUF_X2 inst_16759 ( .A(net_16606), .Z(net_16607) );
DFFR_X2 inst_7131 ( .QN(net_7605), .D(net_3085), .CK(net_9774), .RN(x6501) );
NAND4_X2 inst_3804 ( .ZN(net_3622), .A1(net_3471), .A2(net_3470), .A3(net_3469), .A4(net_3468) );
SDFFR_X2 inst_2266 ( .SI(net_7376), .SE(net_2793), .Q(net_235), .D(net_235), .CK(net_13713), .RN(x6501) );
CLKBUF_X2 inst_17741 ( .A(net_9792), .Z(net_17589) );
CLKBUF_X2 inst_14331 ( .A(net_14178), .Z(net_14179) );
DFFR_X2 inst_7148 ( .QN(net_8948), .D(net_2893), .CK(net_14486), .RN(x6501) );
CLKBUF_X2 inst_13206 ( .A(net_13053), .Z(net_13054) );
CLKBUF_X2 inst_16250 ( .A(net_13712), .Z(net_16098) );
CLKBUF_X2 inst_13440 ( .A(net_13287), .Z(net_13288) );
CLKBUF_X2 inst_15962 ( .A(net_15809), .Z(net_15810) );
AOI221_X2 inst_8744 ( .ZN(net_5658), .B2(net_5657), .C2(net_5655), .A(net_5585), .C1(net_2957), .B1(net_583) );
CLKBUF_X2 inst_12023 ( .A(net_11870), .Z(net_11871) );
CLKBUF_X2 inst_16814 ( .A(net_11852), .Z(net_16662) );
CLKBUF_X2 inst_13437 ( .A(net_13284), .Z(net_13285) );
SDFFR_X2 inst_2514 ( .D(net_7368), .SE(net_2500), .SI(net_232), .Q(net_232), .CK(net_16101), .RN(x6501) );
AOI22_X2 inst_7869 ( .B2(net_4881), .A2(net_4809), .ZN(net_4572), .A1(net_628), .B1(net_234) );
SDFF_X2 inst_1128 ( .D(net_7334), .SI(net_6576), .Q(net_6576), .SE(net_3070), .CK(net_9750) );
AOI22_X2 inst_8009 ( .B1(net_7928), .A1(net_7826), .B2(net_6103), .A2(net_4398), .ZN(net_4126) );
NOR4_X2 inst_3222 ( .ZN(net_2472), .A3(net_2408), .A4(net_2240), .A1(net_1098), .A2(net_1086) );
NAND4_X2 inst_3759 ( .ZN(net_4262), .A1(net_3838), .A2(net_3837), .A3(net_3836), .A4(net_3835) );
CLKBUF_X2 inst_10928 ( .A(net_10775), .Z(net_10776) );
DFFR_X1 inst_7422 ( .QN(net_7506), .D(net_4972), .CK(net_14519), .RN(x6501) );
CLKBUF_X2 inst_19042 ( .A(net_18398), .Z(net_18890) );
NAND2_X2 inst_4070 ( .A2(net_6787), .ZN(net_5777), .A1(net_5775) );
SDFF_X2 inst_1924 ( .D(net_7271), .SI(net_6968), .Q(net_6968), .SE(net_6283), .CK(net_14081) );
CLKBUF_X2 inst_10502 ( .A(net_9171), .Z(net_10350) );
CLKBUF_X2 inst_18452 ( .A(net_18299), .Z(net_18300) );
NAND2_X2 inst_4748 ( .ZN(net_2705), .A2(net_1586), .A1(net_936) );
NAND2_X2 inst_4160 ( .ZN(net_5353), .A1(net_5203), .A2(net_4994) );
INV_X4 inst_5685 ( .A(net_7648), .ZN(net_3082) );
SDFF_X2 inst_961 ( .SI(net_7319), .Q(net_6693), .D(net_6693), .SE(net_3125), .CK(net_9885) );
NOR3_X2 inst_3255 ( .ZN(net_5533), .A3(net_5272), .A1(net_2841), .A2(net_2840) );
CLKBUF_X2 inst_13119 ( .A(net_9295), .Z(net_12967) );
CLKBUF_X2 inst_11082 ( .A(net_10929), .Z(net_10930) );
CLKBUF_X2 inst_12800 ( .A(net_12647), .Z(net_12648) );
AOI22_X2 inst_8077 ( .A1(net_7971), .B1(net_7801), .A2(net_6092), .B2(net_6091), .ZN(net_4067) );
AOI22_X2 inst_8332 ( .B1(net_8883), .A1(net_8328), .B2(net_6252), .A2(net_4345), .ZN(net_3714) );
INV_X4 inst_5103 ( .ZN(net_5683), .A(net_5604) );
CLKBUF_X2 inst_11364 ( .A(net_11211), .Z(net_11212) );
CLKBUF_X2 inst_16734 ( .A(net_15451), .Z(net_16582) );
AOI22_X2 inst_8489 ( .B1(net_6744), .A1(net_6711), .B2(net_6202), .A2(net_3520), .ZN(net_3451) );
SDFFR_X2 inst_2316 ( .SE(net_2260), .Q(net_311), .D(net_311), .CK(net_10467), .RN(x6501), .SI(x3485) );
SDFFR_X1 inst_2737 ( .SI(net_9019), .Q(net_9019), .D(net_7448), .SE(net_3208), .CK(net_10104), .RN(x6501) );
INV_X1 inst_6654 ( .A(net_6151), .ZN(net_6150) );
CLKBUF_X2 inst_14266 ( .A(net_14113), .Z(net_14114) );
SDFF_X2 inst_499 ( .SI(net_8625), .Q(net_8625), .SE(net_3984), .D(net_3950), .CK(net_13268) );
INV_X2 inst_6175 ( .ZN(net_5916), .A(net_5869) );
CLKBUF_X2 inst_9468 ( .A(net_9090), .Z(net_9316) );
SDFFR_X2 inst_2400 ( .SI(net_7370), .SE(net_2732), .D(net_2697), .QN(net_145), .CK(net_16110), .RN(x6501) );
CLKBUF_X2 inst_18535 ( .A(net_18382), .Z(net_18383) );
SDFF_X2 inst_1451 ( .SI(net_7268), .Q(net_7085), .D(net_7085), .SE(net_6278), .CK(net_17076) );
NAND2_X2 inst_4082 ( .A2(net_6761), .A1(net_5835), .ZN(net_5764) );
NAND2_X2 inst_4781 ( .ZN(net_1601), .A2(net_1480), .A1(net_1341) );
CLKBUF_X2 inst_14207 ( .A(net_14054), .Z(net_14055) );
CLKBUF_X2 inst_17779 ( .A(net_17626), .Z(net_17627) );
SDFF_X2 inst_2009 ( .SI(net_7793), .Q(net_7793), .D(net_2713), .SE(net_2459), .CK(net_14243) );
SDFF_X2 inst_501 ( .SI(net_8627), .Q(net_8627), .SE(net_3984), .D(net_3939), .CK(net_10574) );
SDFFS_X2 inst_2093 ( .SI(net_6839), .Q(net_6839), .D(net_6821), .SE(net_2146), .CK(net_18668), .SN(x6501) );
SDFF_X2 inst_1081 ( .D(net_7332), .SI(net_6508), .Q(net_6508), .SE(net_3071), .CK(net_9063) );
OAI211_X2 inst_3195 ( .A(net_7485), .ZN(net_3147), .B(net_3146), .C2(net_2913), .C1(net_2827) );
AOI21_X2 inst_8873 ( .ZN(net_5924), .A(net_5922), .B2(net_5871), .B1(net_2677) );
CLKBUF_X2 inst_10731 ( .A(net_10578), .Z(net_10579) );
CLKBUF_X2 inst_17984 ( .A(net_17831), .Z(net_17832) );
CLKBUF_X2 inst_15888 ( .A(net_15735), .Z(net_15736) );
CLKBUF_X2 inst_15828 ( .A(net_12303), .Z(net_15676) );
OAI33_X1 inst_2905 ( .B2(net_3161), .ZN(net_3019), .B3(net_2912), .A1(net_2850), .B1(net_2773), .A3(net_2591), .A2(net_2531) );
OR2_X4 inst_2819 ( .A2(net_4393), .ZN(net_4392), .A1(net_4391) );
CLKBUF_X2 inst_12263 ( .A(net_12024), .Z(net_12111) );
INV_X2 inst_6293 ( .ZN(net_4205), .A(net_3914) );
CLKBUF_X2 inst_15016 ( .A(net_14863), .Z(net_14864) );
CLKBUF_X2 inst_17416 ( .A(net_17263), .Z(net_17264) );
CLKBUF_X2 inst_9963 ( .A(net_9810), .Z(net_9811) );
SDFF_X2 inst_1114 ( .D(net_7316), .SI(net_6525), .Q(net_6525), .SE(net_3086), .CK(net_12082) );
AOI22_X2 inst_7982 ( .B1(net_8129), .A1(net_7891), .A2(net_6098), .B2(net_4190), .ZN(net_4149) );
CLKBUF_X2 inst_9327 ( .A(net_9138), .Z(net_9175) );
NAND2_X2 inst_4163 ( .ZN(net_5349), .A1(net_5201), .A2(net_4993) );
CLKBUF_X2 inst_15391 ( .A(net_13064), .Z(net_15239) );
AOI211_X2 inst_9020 ( .ZN(net_1918), .B(net_1656), .C2(net_1655), .A(net_1287), .C1(net_1286) );
CLKBUF_X2 inst_17244 ( .A(net_9937), .Z(net_17092) );
CLKBUF_X2 inst_17021 ( .A(net_16073), .Z(net_16869) );
SDFF_X2 inst_1982 ( .D(net_7296), .SI(net_7033), .Q(net_7033), .SE(net_6277), .CK(net_15387) );
CLKBUF_X2 inst_16246 ( .A(net_16093), .Z(net_16094) );
CLKBUF_X2 inst_15909 ( .A(net_11840), .Z(net_15757) );
CLKBUF_X2 inst_11805 ( .A(net_11652), .Z(net_11653) );
SDFF_X2 inst_1849 ( .D(net_7269), .SI(net_6886), .Q(net_6886), .SE(net_6284), .CK(net_16805) );
CLKBUF_X2 inst_18378 ( .A(net_12319), .Z(net_18226) );
INV_X4 inst_5540 ( .ZN(net_1523), .A(net_1106) );
CLKBUF_X2 inst_11123 ( .A(net_10970), .Z(net_10971) );
SDFF_X2 inst_1976 ( .D(net_7272), .SI(net_6849), .Q(net_6849), .SE(net_6282), .CK(net_14069) );
MUX2_X2 inst_4932 ( .A(net_6154), .Z(net_3117), .S(net_2996), .B(net_1207) );
SDFFR_X1 inst_2744 ( .SI(net_9047), .Q(net_9047), .SE(net_3208), .D(net_3113), .CK(net_12932), .RN(x6501) );
NAND4_X2 inst_3681 ( .A4(net_6061), .A1(net_6060), .ZN(net_4584), .A2(net_4004), .A3(net_4003) );
DFFS_X2 inst_6909 ( .QN(net_6804), .D(net_6801), .CK(net_9622), .SN(x6501) );
CLKBUF_X2 inst_13238 ( .A(net_13085), .Z(net_13086) );
INV_X4 inst_5277 ( .ZN(net_1862), .A(net_1773) );
SDFFR_X2 inst_2384 ( .SE(net_2260), .Q(net_321), .D(net_321), .CK(net_10420), .RN(x6501), .SI(x3079) );
NAND2_X2 inst_4614 ( .A2(net_6144), .ZN(net_2613), .A1(net_2612) );
CLKBUF_X2 inst_9606 ( .A(net_9248), .Z(net_9454) );
SDFF_X2 inst_1212 ( .Q(net_7971), .D(net_7971), .SE(net_2755), .SI(net_2660), .CK(net_17038) );
SDFF_X2 inst_670 ( .Q(net_8414), .D(net_8414), .SI(net_3947), .SE(net_3934), .CK(net_12443) );
CLKBUF_X2 inst_17561 ( .A(net_17408), .Z(net_17409) );
NAND2_X2 inst_4180 ( .ZN(net_5324), .A2(net_5190), .A1(net_5075) );
INV_X4 inst_5789 ( .A(net_8262), .ZN(net_2993) );
CLKBUF_X2 inst_11105 ( .A(net_10952), .Z(net_10953) );
CLKBUF_X2 inst_9612 ( .A(net_9369), .Z(net_9460) );
NAND3_X2 inst_3901 ( .ZN(net_5637), .A1(net_5566), .A3(net_5500), .A2(net_5390) );
CLKBUF_X2 inst_18425 ( .A(net_18272), .Z(net_18273) );
CLKBUF_X2 inst_19071 ( .A(net_15367), .Z(net_18919) );
CLKBUF_X2 inst_16901 ( .A(net_16748), .Z(net_16749) );
CLKBUF_X2 inst_17979 ( .A(net_17826), .Z(net_17827) );
HA_X1 inst_6679 ( .S(net_3100), .CO(net_3099), .A(net_3098), .B(net_3087) );
CLKBUF_X2 inst_15200 ( .A(net_15047), .Z(net_15048) );
CLKBUF_X2 inst_14093 ( .A(net_13940), .Z(net_13941) );
INV_X4 inst_5898 ( .A(net_7487), .ZN(net_2935) );
AOI222_X1 inst_8647 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3919), .B1(net_3049), .C1(net_3048), .A1(x13786) );
CLKBUF_X2 inst_10845 ( .A(net_9632), .Z(net_10693) );
CLKBUF_X2 inst_9814 ( .A(net_9370), .Z(net_9662) );
CLKBUF_X2 inst_14502 ( .A(net_11546), .Z(net_14350) );
SDFF_X2 inst_807 ( .SI(net_8496), .Q(net_8496), .D(net_3959), .SE(net_3884), .CK(net_9983) );
SDFF_X2 inst_705 ( .SI(net_8598), .Q(net_8598), .SE(net_3984), .D(net_3965), .CK(net_13033) );
CLKBUF_X2 inst_18433 ( .A(net_18280), .Z(net_18281) );
SDFF_X2 inst_911 ( .SI(net_8730), .Q(net_8730), .SE(net_6195), .D(net_3975), .CK(net_10215) );
CLKBUF_X2 inst_10921 ( .A(net_10768), .Z(net_10769) );
CLKBUF_X2 inst_15746 ( .A(net_12912), .Z(net_15594) );
SDFF_X2 inst_1003 ( .D(net_7310), .SI(net_6651), .Q(net_6651), .SE(net_3123), .CK(net_11906) );
CLKBUF_X2 inst_14893 ( .A(net_14740), .Z(net_14741) );
CLKBUF_X2 inst_13804 ( .A(net_13651), .Z(net_13652) );
CLKBUF_X2 inst_14889 ( .A(net_14736), .Z(net_14737) );
CLKBUF_X2 inst_10284 ( .A(net_9413), .Z(net_10132) );
NOR2_X2 inst_3469 ( .ZN(net_2553), .A2(net_2496), .A1(net_2454) );
INV_X4 inst_6026 ( .A(net_6313), .ZN(net_2679) );
INV_X4 inst_5456 ( .ZN(net_852), .A(net_777) );
SDFFS_X2 inst_2080 ( .SI(net_7378), .SE(net_2794), .Q(net_167), .D(net_167), .CK(net_13668), .SN(x6501) );
SDFF_X2 inst_1625 ( .Q(net_8168), .D(net_8168), .SI(net_2712), .SE(net_2538), .CK(net_13771) );
SDFF_X2 inst_593 ( .SI(net_8385), .Q(net_8385), .SE(net_3969), .D(net_3959), .CK(net_10161) );
INV_X4 inst_5707 ( .ZN(net_2547), .A(net_260) );
CLKBUF_X2 inst_18920 ( .A(net_18517), .Z(net_18768) );
CLKBUF_X2 inst_15664 ( .A(net_15511), .Z(net_15512) );
SDFFR_X2 inst_2223 ( .Q(net_7452), .D(net_7452), .SE(net_2863), .CK(net_12918), .SI(x13560), .RN(x6501) );
NAND2_X2 inst_4522 ( .ZN(net_3569), .A2(net_3568), .A1(net_3561) );
INV_X4 inst_6137 ( .A(net_6113), .ZN(net_6111) );
CLKBUF_X2 inst_12426 ( .A(net_12273), .Z(net_12274) );
CLKBUF_X2 inst_10099 ( .A(net_9946), .Z(net_9947) );
INV_X4 inst_5738 ( .A(net_7374), .ZN(net_931) );
AOI22_X2 inst_7845 ( .A2(net_5595), .ZN(net_4663), .B2(net_4388), .B1(net_2630), .A1(net_314) );
AND2_X4 inst_9065 ( .ZN(net_6202), .A2(net_3250), .A1(net_3249) );
CLKBUF_X2 inst_10045 ( .A(net_9892), .Z(net_9893) );
SDFF_X2 inst_479 ( .SI(net_8453), .Q(net_8453), .SE(net_3983), .D(net_3937), .CK(net_11102) );
CLKBUF_X2 inst_10448 ( .A(net_10295), .Z(net_10296) );
CLKBUF_X2 inst_17271 ( .A(net_17118), .Z(net_17119) );
SDFFR_X2 inst_2344 ( .D(net_7366), .SE(net_2734), .SI(net_272), .Q(net_272), .CK(net_13689), .RN(x6501) );
NOR2_X4 inst_3326 ( .ZN(net_3381), .A2(net_3260), .A1(net_3259) );
DFFR_X2 inst_7288 ( .Q(net_7301), .D(net_1683), .CK(net_18717), .RN(x6501) );
CLKBUF_X2 inst_12892 ( .A(net_9172), .Z(net_12740) );
NAND2_X2 inst_4387 ( .A1(net_7119), .A2(net_5164), .ZN(net_5070) );
CLKBUF_X2 inst_9420 ( .A(net_9267), .Z(net_9268) );
CLKBUF_X2 inst_15068 ( .A(net_14915), .Z(net_14916) );
DFFR_X2 inst_7113 ( .QN(net_7611), .D(net_3094), .CK(net_11226), .RN(x6501) );
INV_X4 inst_5780 ( .A(net_7588), .ZN(net_551) );
CLKBUF_X2 inst_16485 ( .A(net_10867), .Z(net_16333) );
CLKBUF_X2 inst_10523 ( .A(net_10370), .Z(net_10371) );
CLKBUF_X2 inst_17320 ( .A(net_17167), .Z(net_17168) );
NAND2_X2 inst_4497 ( .ZN(net_4473), .A2(net_4468), .A1(net_1801) );
SDFFR_X1 inst_2651 ( .D(net_6774), .SE(net_4506), .CK(net_9197), .RN(x6501), .SI(x1667), .Q(x1667) );
NAND2_X2 inst_4756 ( .A2(net_2204), .ZN(net_1754), .A1(net_1537) );
NAND2_X2 inst_4201 ( .ZN(net_5296), .A2(net_5176), .A1(net_5054) );
INV_X4 inst_5658 ( .A(net_7370), .ZN(net_1122) );
XOR2_X2 inst_48 ( .B(net_3145), .A(net_1457), .Z(net_1014) );
CLKBUF_X2 inst_16008 ( .A(net_15855), .Z(net_15856) );
SDFFR_X2 inst_2246 ( .SI(net_7374), .SE(net_2793), .Q(net_233), .D(net_233), .CK(net_13717), .RN(x6501) );
DFFR_X1 inst_7507 ( .D(net_1888), .Q(net_258), .CK(net_14846), .RN(x6501) );
SDFF_X2 inst_443 ( .Q(net_8772), .D(net_8772), .SE(net_3982), .SI(net_3951), .CK(net_13435) );
CLKBUF_X2 inst_17114 ( .A(net_13488), .Z(net_16962) );
CLKBUF_X2 inst_11022 ( .A(net_10869), .Z(net_10870) );
AOI221_X2 inst_8766 ( .C1(net_8988), .B2(net_5538), .ZN(net_5457), .C2(net_5456), .A(net_4944), .B1(net_417) );
NAND2_X2 inst_4259 ( .A1(net_6911), .A2(net_5247), .ZN(net_5201) );
CLKBUF_X2 inst_12152 ( .A(net_11999), .Z(net_12000) );
AND2_X4 inst_9060 ( .A1(net_3328), .ZN(net_3306), .A2(net_3305) );
SDFF_X2 inst_1700 ( .Q(net_8189), .D(net_8189), .SI(net_2573), .SE(net_2561), .CK(net_15260) );
CLKBUF_X2 inst_15814 ( .A(net_12802), .Z(net_15662) );
SDFFR_X2 inst_2571 ( .SI(net_6832), .Q(net_6832), .D(net_6829), .SE(net_2146), .CK(net_18690), .RN(x6501) );
CLKBUF_X2 inst_12481 ( .A(net_12328), .Z(net_12329) );
SDFF_X2 inst_730 ( .SI(net_8366), .Q(net_8366), .D(net_3950), .SE(net_3880), .CK(net_10532) );
CLKBUF_X2 inst_11430 ( .A(net_11277), .Z(net_11278) );
CLKBUF_X2 inst_10116 ( .A(net_9963), .Z(net_9964) );
DFF_X1 inst_6754 ( .Q(net_6764), .D(net_5612), .CK(net_11542) );
XNOR2_X2 inst_321 ( .A(net_1779), .ZN(net_940), .B(net_939) );
CLKBUF_X2 inst_18831 ( .A(net_18678), .Z(net_18679) );
CLKBUF_X2 inst_10977 ( .A(net_9399), .Z(net_10825) );
CLKBUF_X2 inst_18085 ( .A(net_17932), .Z(net_17933) );
OAI21_X2 inst_3131 ( .ZN(net_2388), .A(net_2179), .B2(net_2161), .B1(net_1639) );
CLKBUF_X2 inst_12684 ( .A(net_9077), .Z(net_12532) );
CLKBUF_X2 inst_14788 ( .A(net_14635), .Z(net_14636) );
CLKBUF_X2 inst_13308 ( .A(net_12090), .Z(net_13156) );
AOI22_X2 inst_8264 ( .A1(net_8616), .B1(net_8431), .A2(net_3864), .B2(net_3863), .ZN(net_3774) );
CLKBUF_X2 inst_16049 ( .A(net_14277), .Z(net_15897) );
CLKBUF_X2 inst_16834 ( .A(net_11446), .Z(net_16682) );
SDFF_X2 inst_1152 ( .SI(net_7333), .Q(net_6608), .D(net_6608), .SE(net_3069), .CK(net_11671) );
DFFS_X2 inst_6878 ( .Q(net_6460), .D(net_3338), .CK(net_15084), .SN(x6501) );
CLKBUF_X2 inst_15255 ( .A(net_15102), .Z(net_15103) );
INV_X2 inst_6517 ( .ZN(net_814), .A(net_219) );
CLKBUF_X2 inst_18582 ( .A(net_18429), .Z(net_18430) );
DFF_X1 inst_6823 ( .QN(net_8237), .D(net_4444), .CK(net_17198) );
AOI222_X1 inst_8670 ( .C2(net_5832), .A2(net_5830), .B2(net_5824), .ZN(net_3585), .A1(net_3266), .B1(net_2148), .C1(x2542) );
XNOR2_X2 inst_182 ( .ZN(net_1672), .B(net_1581), .A(net_1580) );
SDFF_X2 inst_931 ( .SI(net_8704), .Q(net_8704), .SE(net_6195), .D(net_3961), .CK(net_10122) );
AND2_X2 inst_9205 ( .ZN(net_2540), .A1(net_510), .A2(net_497) );
OAI21_X1 inst_3174 ( .B2(net_4221), .ZN(net_3971), .A(net_3230), .B1(net_3187) );
SDFF_X2 inst_1674 ( .SI(net_7743), .Q(net_7743), .D(net_2659), .SE(net_2560), .CK(net_18534) );
NAND4_X2 inst_3824 ( .ZN(net_3047), .A4(net_3046), .A3(net_3038), .A1(x2355), .A2(x2308) );
DFFS_X2 inst_6895 ( .Q(net_6319), .D(net_2636), .CK(net_17460), .SN(x6501) );
CLKBUF_X2 inst_12807 ( .A(net_12654), .Z(net_12655) );
AOI22_X2 inst_8438 ( .B1(net_6666), .A1(net_6633), .A2(net_6213), .B2(net_6138), .ZN(net_3503) );
CLKBUF_X2 inst_15983 ( .A(net_15830), .Z(net_15831) );
AOI22_X2 inst_8315 ( .B1(net_8780), .A1(net_8521), .A2(net_3861), .B2(net_3860), .ZN(net_3730) );
CLKBUF_X2 inst_16226 ( .A(net_16073), .Z(net_16074) );
NAND2_X2 inst_4089 ( .ZN(net_5450), .A1(net_5170), .A2(net_5169) );
CLKBUF_X2 inst_15929 ( .A(net_15776), .Z(net_15777) );
CLKBUF_X2 inst_14320 ( .A(net_10316), .Z(net_14168) );
SDFF_X2 inst_1415 ( .Q(net_7156), .D(net_7156), .SE(net_6279), .SI(net_2544), .CK(net_15901) );
CLKBUF_X2 inst_12089 ( .A(net_11936), .Z(net_11937) );
CLKBUF_X2 inst_13631 ( .A(net_13478), .Z(net_13479) );
NOR3_X2 inst_3301 ( .A3(net_2733), .ZN(net_1818), .A2(net_1817), .A1(net_1660) );
INV_X4 inst_5997 ( .A(net_7665), .ZN(net_1643) );
INV_X2 inst_6469 ( .A(net_7587), .ZN(net_3136) );
CLKBUF_X2 inst_12571 ( .A(net_12418), .Z(net_12419) );
CLKBUF_X2 inst_19164 ( .A(net_11336), .Z(net_19012) );
CLKBUF_X2 inst_13433 ( .A(net_11730), .Z(net_13281) );
INV_X4 inst_5578 ( .A(net_6375), .ZN(net_617) );
CLKBUF_X2 inst_13396 ( .A(net_13243), .Z(net_13244) );
AOI222_X1 inst_8655 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3911), .B1(net_1674), .C1(net_1673), .A1(x13884) );
CLKBUF_X2 inst_11459 ( .A(net_10815), .Z(net_11307) );
NAND2_X2 inst_4599 ( .A2(net_2943), .ZN(net_2772), .A1(net_2652) );
AOI22_X2 inst_8147 ( .B1(net_8052), .A1(net_7848), .B2(net_6107), .ZN(net_6061), .A2(net_4400) );
INV_X4 inst_5906 ( .ZN(net_2501), .A(net_339) );
NAND2_X2 inst_4677 ( .A1(net_9008), .A2(net_6164), .ZN(net_2264) );
CLKBUF_X2 inst_14796 ( .A(net_12222), .Z(net_14644) );
INV_X4 inst_5516 ( .ZN(net_862), .A(net_677) );
SDFF_X2 inst_1698 ( .SI(net_7290), .Q(net_7067), .D(net_7067), .SE(net_6280), .CK(net_18264) );
CLKBUF_X2 inst_11698 ( .A(net_11545), .Z(net_11546) );
SDFF_X2 inst_944 ( .SI(net_7326), .Q(net_6700), .D(net_6700), .SE(net_3125), .CK(net_11304) );
INV_X4 inst_5248 ( .ZN(net_2161), .A(net_1869) );
CLKBUF_X2 inst_15488 ( .A(net_10421), .Z(net_15336) );
AOI22_X2 inst_7992 ( .B1(net_8028), .A1(net_7994), .B2(net_6102), .A2(net_6097), .ZN(net_4140) );
CLKBUF_X2 inst_16924 ( .A(net_12411), .Z(net_16772) );
SDFF_X2 inst_459 ( .SI(net_8462), .Q(net_8462), .SE(net_3983), .D(net_3967), .CK(net_10187) );
AOI22_X2 inst_8259 ( .B1(net_8800), .A1(net_8541), .A2(net_3861), .B2(net_3860), .ZN(net_3779) );
CLKBUF_X2 inst_11737 ( .A(net_11584), .Z(net_11585) );
AOI22_X2 inst_8532 ( .B1(net_6525), .A1(net_6492), .A2(net_6137), .B2(net_6104), .ZN(net_3408) );
CLKBUF_X2 inst_10084 ( .A(net_9931), .Z(net_9932) );
DFFR_X1 inst_7461 ( .D(net_4680), .CK(net_9590), .RN(x6501), .Q(x1107) );
CLKBUF_X2 inst_12861 ( .A(net_11009), .Z(net_12709) );
CLKBUF_X2 inst_17396 ( .A(net_17243), .Z(net_17244) );
CLKBUF_X2 inst_13723 ( .A(net_10353), .Z(net_13571) );
NOR2_X2 inst_3393 ( .ZN(net_4905), .A2(net_4411), .A1(net_4408) );
AOI222_X1 inst_8613 ( .B2(net_6759), .B1(net_5835), .A2(net_5830), .C2(net_5824), .ZN(net_5800), .C1(net_2128), .A1(net_1313) );
CLKBUF_X2 inst_18470 ( .A(net_10907), .Z(net_18318) );
AOI22_X2 inst_8148 ( .A1(net_7950), .B1(net_7780), .A2(net_6092), .B2(net_6091), .ZN(net_4004) );
CLKBUF_X2 inst_18403 ( .A(net_18250), .Z(net_18251) );
MUX2_X2 inst_4976 ( .A(net_9045), .B(net_7442), .Z(net_3940), .S(net_622) );
CLKBUF_X2 inst_9657 ( .A(net_9123), .Z(net_9505) );
NOR2_X2 inst_3409 ( .A1(net_6256), .ZN(net_3566), .A2(net_3304) );
CLKBUF_X2 inst_13252 ( .A(net_11812), .Z(net_13100) );
NOR2_X2 inst_3591 ( .A1(net_7353), .A2(net_1446), .ZN(net_1164) );
INV_X4 inst_5970 ( .A(net_6754), .ZN(net_1508) );
CLKBUF_X2 inst_16888 ( .A(net_16735), .Z(net_16736) );
CLKBUF_X2 inst_16242 ( .A(net_16076), .Z(net_16090) );
SDFF_X2 inst_450 ( .Q(net_8747), .D(net_8747), .SE(net_3982), .SI(net_3947), .CK(net_12475) );
CLKBUF_X2 inst_9723 ( .A(net_9131), .Z(net_9571) );
CLKBUF_X2 inst_18785 ( .A(net_18632), .Z(net_18633) );
SDFF_X2 inst_520 ( .Q(net_8874), .D(net_8874), .SI(net_3963), .SE(net_3936), .CK(net_10077) );
INV_X4 inst_5717 ( .A(net_8914), .ZN(net_4666) );
NAND4_X2 inst_3658 ( .A4(net_6008), .A1(net_6007), .ZN(net_4607), .A2(net_4144), .A3(net_4143) );
CLKBUF_X2 inst_10019 ( .A(net_9866), .Z(net_9867) );
CLKBUF_X2 inst_18701 ( .A(net_18548), .Z(net_18549) );
CLKBUF_X2 inst_17142 ( .A(net_9319), .Z(net_16990) );
CLKBUF_X2 inst_11667 ( .A(net_9227), .Z(net_11515) );
NAND2_X2 inst_4554 ( .A1(net_7513), .ZN(net_3276), .A2(net_3263) );
CLKBUF_X2 inst_14850 ( .A(net_14697), .Z(net_14698) );
INV_X4 inst_5977 ( .A(net_7233), .ZN(net_1856) );
SDFF_X2 inst_2026 ( .SI(net_7941), .Q(net_7941), .D(net_2703), .SE(net_2461), .CK(net_16702) );
NAND4_X4 inst_3623 ( .ZN(net_6158), .A4(net_5983), .A1(net_5982), .A3(net_2410), .A2(net_2173) );
SDFF_X2 inst_1556 ( .Q(net_7985), .D(net_7985), .SI(net_2573), .SE(net_2542), .CK(net_15273) );
CLKBUF_X2 inst_9228 ( .A(net_9075), .Z(net_9076) );
CLKBUF_X2 inst_14820 ( .A(net_14667), .Z(net_14668) );
DFF_X1 inst_6796 ( .QN(net_8243), .D(net_4437), .CK(net_17596) );
CLKBUF_X2 inst_15636 ( .A(net_15483), .Z(net_15484) );
CLKBUF_X2 inst_11243 ( .A(net_11090), .Z(net_11091) );
CLKBUF_X2 inst_17450 ( .A(net_17297), .Z(net_17298) );
CLKBUF_X2 inst_12075 ( .A(net_11922), .Z(net_11923) );
CLKBUF_X2 inst_14410 ( .A(net_11962), .Z(net_14258) );
SDFF_X2 inst_862 ( .Q(net_8570), .D(net_8570), .SI(net_3959), .SE(net_3878), .CK(net_13163) );
NAND2_X2 inst_4358 ( .A1(net_7042), .A2(net_5162), .ZN(net_5099) );
NAND2_X2 inst_4390 ( .A1(net_7083), .A2(net_5164), .ZN(net_5067) );
CLKBUF_X2 inst_16387 ( .A(net_16234), .Z(net_16235) );
CLKBUF_X2 inst_14618 ( .A(net_14465), .Z(net_14466) );
CLKBUF_X2 inst_17383 ( .A(net_17230), .Z(net_17231) );
CLKBUF_X2 inst_10620 ( .A(net_9364), .Z(net_10468) );
SDFF_X2 inst_1764 ( .SI(net_8048), .Q(net_8048), .D(net_2709), .SE(net_2508), .CK(net_15734) );
CLKBUF_X2 inst_14024 ( .A(net_13871), .Z(net_13872) );
INV_X4 inst_5271 ( .A(net_1861), .ZN(net_1691) );
CLKBUF_X2 inst_14799 ( .A(net_14646), .Z(net_14647) );
INV_X4 inst_5323 ( .A(net_2652), .ZN(net_2307) );
CLKBUF_X2 inst_15366 ( .A(net_15213), .Z(net_15214) );
DFFR_X1 inst_7472 ( .QN(net_7425), .D(net_4023), .CK(net_12395), .RN(x6501) );
SDFF_X2 inst_1159 ( .SI(net_7342), .Q(net_6617), .D(net_6617), .SE(net_3069), .CK(net_11666) );
AOI221_X2 inst_8740 ( .ZN(net_5749), .B2(net_5657), .A(net_5611), .C2(net_5535), .B1(net_2698), .C1(net_446) );
CLKBUF_X2 inst_9550 ( .A(net_9215), .Z(net_9398) );
AOI222_X1 inst_8659 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3907), .B1(net_3331), .C1(net_3330), .A1(x13808) );
CLKBUF_X2 inst_16612 ( .A(net_16459), .Z(net_16460) );
CLKBUF_X2 inst_9835 ( .A(net_9682), .Z(net_9683) );
SDFF_X2 inst_938 ( .SI(net_7316), .Q(net_6657), .D(net_6657), .SE(net_3126), .CK(net_12155) );
CLKBUF_X2 inst_16420 ( .A(net_10266), .Z(net_16268) );
CLKBUF_X2 inst_14521 ( .A(net_12415), .Z(net_14369) );
CLKBUF_X2 inst_11189 ( .A(net_9188), .Z(net_11037) );
CLKBUF_X2 inst_12552 ( .A(net_12399), .Z(net_12400) );
CLKBUF_X2 inst_12742 ( .A(net_12589), .Z(net_12590) );
CLKBUF_X2 inst_16752 ( .A(net_12412), .Z(net_16600) );
INV_X16 inst_6646 ( .ZN(net_6098), .A(net_3569) );
CLKBUF_X2 inst_9698 ( .A(net_9117), .Z(net_9546) );
NAND4_X2 inst_3638 ( .ZN(net_5026), .A4(net_4770), .A1(net_4700), .A3(net_4687), .A2(net_4670) );
AOI21_X2 inst_8923 ( .B2(net_5871), .ZN(net_5701), .A(net_5700), .B1(x577) );
NAND2_X2 inst_4365 ( .A1(net_7152), .A2(net_5166), .ZN(net_5092) );
CLKBUF_X2 inst_9399 ( .A(net_9246), .Z(net_9247) );
CLKBUF_X2 inst_18899 ( .A(net_18746), .Z(net_18747) );
CLKBUF_X2 inst_16881 ( .A(net_16728), .Z(net_16729) );
CLKBUF_X2 inst_18151 ( .A(net_17998), .Z(net_17999) );
AOI21_X2 inst_8957 ( .B2(net_5609), .ZN(net_5274), .A(net_4941), .B1(net_377) );
CLKBUF_X2 inst_11320 ( .A(net_11124), .Z(net_11168) );
CLKBUF_X2 inst_14253 ( .A(net_14100), .Z(net_14101) );
CLKBUF_X2 inst_19124 ( .A(net_18971), .Z(net_18972) );
DFFR_X1 inst_7426 ( .QN(net_8927), .D(net_4861), .CK(net_17328), .RN(x6501) );
SDFFS_X1 inst_2102 ( .D(net_9054), .SI(net_7594), .Q(net_7594), .SE(net_3144), .CK(net_13444), .SN(x6501) );
CLKBUF_X2 inst_14070 ( .A(net_13917), .Z(net_13918) );
CLKBUF_X2 inst_9762 ( .A(net_9424), .Z(net_9610) );
NAND2_X2 inst_4908 ( .A2(net_7376), .ZN(net_603), .A1(net_165) );
DFFR_X2 inst_7160 ( .QN(net_7221), .D(net_2766), .CK(net_18952), .RN(x6501) );
CLKBUF_X2 inst_10343 ( .A(net_10190), .Z(net_10191) );
CLKBUF_X2 inst_16806 ( .A(net_16653), .Z(net_16654) );
INV_X32 inst_6168 ( .ZN(net_5162), .A(net_4817) );
AOI22_X2 inst_8445 ( .B1(net_6734), .A1(net_6701), .B2(net_6202), .A2(net_3520), .ZN(net_3495) );
CLKBUF_X2 inst_18892 ( .A(net_18127), .Z(net_18740) );
CLKBUF_X2 inst_11182 ( .A(net_11029), .Z(net_11030) );
SDFF_X2 inst_784 ( .SI(net_8335), .Q(net_8335), .D(net_3943), .SE(net_3880), .CK(net_12948) );
NOR4_X2 inst_3237 ( .ZN(net_1796), .A2(net_1493), .A1(net_1490), .A4(net_812), .A3(net_785) );
SDFF_X2 inst_1264 ( .Q(net_8109), .D(net_8109), .SI(net_2716), .SE(net_2707), .CK(net_17101) );
CLKBUF_X2 inst_19185 ( .A(net_19032), .Z(net_19033) );
SDFF_X2 inst_690 ( .Q(net_8882), .D(net_8882), .SI(net_3940), .SE(net_3936), .CK(net_10247) );
CLKBUF_X2 inst_18469 ( .A(net_18316), .Z(net_18317) );
CLKBUF_X2 inst_11895 ( .A(net_11742), .Z(net_11743) );
SDFF_X2 inst_2025 ( .SI(net_7939), .Q(net_7939), .D(net_2716), .SE(net_2461), .CK(net_16963) );
AOI22_X2 inst_7819 ( .A2(net_8252), .B1(net_5033), .ZN(net_4731), .A1(net_4729), .B2(net_4728) );
CLKBUF_X2 inst_10607 ( .A(net_9528), .Z(net_10455) );
NAND2_X2 inst_4717 ( .ZN(net_6172), .A2(net_6122), .A1(net_1716) );
CLKBUF_X2 inst_12722 ( .A(net_12569), .Z(net_12570) );
CLKBUF_X2 inst_18179 ( .A(net_18026), .Z(net_18027) );
CLKBUF_X2 inst_10969 ( .A(net_10511), .Z(net_10817) );
CLKBUF_X2 inst_9666 ( .A(net_9489), .Z(net_9514) );
XOR2_X1 inst_75 ( .B(net_7516), .Z(net_6177), .A(net_3198) );
CLKBUF_X2 inst_15656 ( .A(net_15503), .Z(net_15504) );
INV_X2 inst_6386 ( .ZN(net_1319), .A(net_1318) );
CLKBUF_X2 inst_16182 ( .A(net_16029), .Z(net_16030) );
AOI22_X2 inst_7986 ( .A1(net_7959), .B1(net_7789), .A2(net_6092), .B2(net_6091), .ZN(net_4145) );
CLKBUF_X2 inst_19046 ( .A(net_18893), .Z(net_18894) );
CLKBUF_X2 inst_9286 ( .A(net_9114), .Z(net_9134) );
AOI22_X2 inst_7891 ( .B1(net_9001), .A2(net_5538), .B2(net_5456), .ZN(net_4539), .A1(net_430) );
CLKBUF_X2 inst_18984 ( .A(net_18831), .Z(net_18832) );
CLKBUF_X2 inst_12082 ( .A(net_11929), .Z(net_11930) );
CLKBUF_X2 inst_19171 ( .A(net_19018), .Z(net_19019) );
CLKBUF_X2 inst_13938 ( .A(net_13785), .Z(net_13786) );
CLKBUF_X2 inst_10890 ( .A(net_10180), .Z(net_10738) );
CLKBUF_X2 inst_10339 ( .A(net_10186), .Z(net_10187) );
SDFF_X2 inst_1024 ( .SI(net_7315), .Q(net_6722), .D(net_6722), .SE(net_3124), .CK(net_12110) );
INV_X4 inst_5827 ( .A(net_7573), .ZN(net_540) );
CLKBUF_X2 inst_12144 ( .A(net_11991), .Z(net_11992) );
SDFFR_X2 inst_2232 ( .Q(net_7466), .D(net_7466), .SE(net_2863), .CK(net_12164), .SI(x13464), .RN(x6501) );
NAND2_X2 inst_4546 ( .ZN(net_3324), .A1(net_3323), .A2(net_3322) );
CLKBUF_X2 inst_13218 ( .A(net_10913), .Z(net_13066) );
CLKBUF_X2 inst_12061 ( .A(net_9401), .Z(net_11909) );
CLKBUF_X2 inst_16716 ( .A(net_16563), .Z(net_16564) );
SDFF_X2 inst_1689 ( .Q(net_8028), .D(net_8028), .SI(net_2590), .SE(net_2545), .CK(net_15582) );
AOI22_X2 inst_8279 ( .A1(net_8618), .B1(net_8433), .A2(net_3864), .B2(net_3863), .ZN(net_3762) );
OR2_X4 inst_2846 ( .ZN(net_4390), .A2(net_1636), .A1(net_1633) );
NOR2_X2 inst_3584 ( .A1(net_8962), .ZN(net_1178), .A2(net_1061) );
CLKBUF_X2 inst_11408 ( .A(net_11255), .Z(net_11256) );
CLKBUF_X2 inst_9472 ( .A(net_9319), .Z(net_9320) );
SDFF_X2 inst_1448 ( .SI(net_7297), .Q(net_7114), .D(net_7114), .SE(net_6278), .CK(net_18205) );
AOI22_X2 inst_8395 ( .A1(net_8599), .B1(net_8414), .A2(net_3864), .B2(net_3863), .ZN(net_3656) );
SDFF_X2 inst_1816 ( .D(net_7267), .SI(net_6924), .Q(net_6924), .SE(net_6281), .CK(net_14128) );
CLKBUF_X2 inst_11892 ( .A(net_11433), .Z(net_11740) );
CLKBUF_X2 inst_11723 ( .A(net_11570), .Z(net_11571) );
CLKBUF_X2 inst_14829 ( .A(net_14676), .Z(net_14677) );
INV_X8 inst_5012 ( .ZN(net_5595), .A(net_4410) );
NOR2_X2 inst_3381 ( .ZN(net_5544), .A1(net_5301), .A2(net_5300) );
CLKBUF_X2 inst_17636 ( .A(net_17483), .Z(net_17484) );
CLKBUF_X2 inst_14123 ( .A(net_13970), .Z(net_13971) );
SDFF_X2 inst_1091 ( .D(net_7316), .SI(net_6492), .Q(net_6492), .SE(net_3071), .CK(net_12087) );
CLKBUF_X2 inst_9915 ( .A(net_9762), .Z(net_9763) );
NAND2_X2 inst_4837 ( .A2(net_7397), .ZN(net_921), .A1(net_908) );
INV_X8 inst_5059 ( .ZN(net_6265), .A(net_3375) );
AOI22_X2 inst_8206 ( .B1(net_8571), .A1(net_8460), .A2(net_6263), .B2(net_6262), .ZN(net_3830) );
CLKBUF_X2 inst_10450 ( .A(net_10297), .Z(net_10298) );
CLKBUF_X2 inst_16308 ( .A(net_16155), .Z(net_16156) );
CLKBUF_X2 inst_13800 ( .A(net_13647), .Z(net_13648) );
CLKBUF_X2 inst_18525 ( .A(net_18372), .Z(net_18373) );
NAND2_X2 inst_4154 ( .ZN(net_5361), .A1(net_5207), .A2(net_4996) );
CLKBUF_X2 inst_10374 ( .A(net_10221), .Z(net_10222) );
INV_X4 inst_5398 ( .A(net_1337), .ZN(net_884) );
NAND2_X2 inst_4816 ( .ZN(net_1248), .A1(net_901), .A2(net_843) );
OAI211_X2 inst_3179 ( .ZN(net_5748), .A(net_5747), .B(net_5598), .C2(net_2947), .C1(net_2912) );
OAI21_X2 inst_3059 ( .B2(net_8243), .B1(net_4850), .ZN(net_4748), .A(net_2633) );
CLKBUF_X2 inst_15297 ( .A(net_12306), .Z(net_15145) );
CLKBUF_X2 inst_11357 ( .A(net_11204), .Z(net_11205) );
CLKBUF_X2 inst_15660 ( .A(net_15507), .Z(net_15508) );
CLKBUF_X2 inst_9390 ( .A(net_9173), .Z(net_9238) );
SDFFR_X2 inst_2587 ( .D(net_7382), .QN(net_7242), .SI(net_1950), .SE(net_1379), .CK(net_14745), .RN(x6501) );
HA_X1 inst_6680 ( .A(net_3239), .S(net_3097), .CO(net_3096), .B(net_2972) );
AOI21_X4 inst_8868 ( .B2(net_6173), .ZN(net_6171), .B1(net_2642), .A(net_1804) );
CLKBUF_X2 inst_13072 ( .A(net_12919), .Z(net_12920) );
AOI21_X2 inst_8883 ( .ZN(net_5845), .A(net_5844), .B2(net_5843), .B1(net_2679) );
OAI21_X2 inst_3031 ( .B1(net_4954), .ZN(net_4930), .B2(net_4847), .A(net_4716) );
CLKBUF_X2 inst_18218 ( .A(net_18065), .Z(net_18066) );
SDFF_X2 inst_1257 ( .Q(net_8091), .D(net_8091), .SI(net_2720), .SE(net_2707), .CK(net_18420) );
SDFF_X2 inst_875 ( .Q(net_8586), .D(net_8586), .SI(net_3940), .SE(net_3878), .CK(net_10220) );
NOR3_X2 inst_3298 ( .ZN(net_2115), .A1(net_1876), .A3(net_1785), .A2(net_1597) );
NOR2_X2 inst_3482 ( .A1(net_2652), .ZN(net_2238), .A2(net_2059) );
INV_X4 inst_5075 ( .ZN(net_5850), .A(net_5797) );
CLKBUF_X2 inst_17680 ( .A(net_17527), .Z(net_17528) );
SDFFS_X2 inst_2069 ( .SI(net_2803), .SE(net_2795), .Q(net_175), .D(net_175), .CK(net_14670), .SN(x6501) );
CLKBUF_X2 inst_15032 ( .A(net_14879), .Z(net_14880) );
NAND2_X2 inst_4098 ( .ZN(net_5436), .A1(net_5158), .A2(net_5157) );
CLKBUF_X2 inst_11220 ( .A(net_11067), .Z(net_11068) );
INV_X4 inst_5703 ( .A(net_8943), .ZN(net_1273) );
OAI21_X4 inst_2978 ( .ZN(net_6187), .B2(net_4512), .A(net_4467), .B1(net_4371) );
CLKBUF_X2 inst_14817 ( .A(net_10771), .Z(net_14665) );
CLKBUF_X2 inst_14239 ( .A(net_14086), .Z(net_14087) );
CLKBUF_X2 inst_11033 ( .A(net_10880), .Z(net_10881) );
CLKBUF_X2 inst_11393 ( .A(net_11164), .Z(net_11241) );
CLKBUF_X2 inst_10269 ( .A(net_10116), .Z(net_10117) );
CLKBUF_X2 inst_14352 ( .A(net_14199), .Z(net_14200) );
SDFF_X2 inst_2019 ( .SI(net_7781), .Q(net_7781), .D(net_2573), .SE(net_2459), .CK(net_18020) );
CLKBUF_X2 inst_13679 ( .A(net_13526), .Z(net_13527) );
AOI22_X2 inst_8323 ( .B1(net_8771), .A1(net_8401), .A2(net_3867), .B2(net_3866), .ZN(net_3723) );
INV_X4 inst_5186 ( .ZN(net_4971), .A(net_4888) );
CLKBUF_X2 inst_15061 ( .A(net_14908), .Z(net_14909) );
XOR2_X1 inst_69 ( .Z(net_3922), .B(net_3921), .A(net_3531) );
CLKBUF_X2 inst_18854 ( .A(net_18701), .Z(net_18702) );
CLKBUF_X2 inst_18077 ( .A(net_17924), .Z(net_17925) );
CLKBUF_X2 inst_15542 ( .A(net_15389), .Z(net_15390) );
CLKBUF_X2 inst_14448 ( .A(net_14295), .Z(net_14296) );
SDFFR_X1 inst_2669 ( .D(net_6786), .SE(net_4506), .CK(net_9179), .RN(x6501), .SI(x1244), .Q(x1244) );
CLKBUF_X2 inst_15396 ( .A(net_15243), .Z(net_15244) );
CLKBUF_X2 inst_17278 ( .A(net_13877), .Z(net_17126) );
CLKBUF_X2 inst_12844 ( .A(net_11762), .Z(net_12692) );
CLKBUF_X2 inst_17319 ( .A(net_11445), .Z(net_17167) );
SDFF_X2 inst_844 ( .SI(net_8656), .Q(net_8656), .D(net_3975), .SE(net_3885), .CK(net_12507) );
SDFFR_X2 inst_2489 ( .Q(net_8972), .D(net_8972), .SI(net_4528), .SE(net_2562), .CK(net_14803), .RN(x6501) );
CLKBUF_X2 inst_14712 ( .A(net_14559), .Z(net_14560) );
DFFR_X2 inst_6968 ( .QN(net_6287), .D(net_5932), .CK(net_13889), .RN(x6501) );
NOR2_X1 inst_3619 ( .A1(net_6163), .ZN(net_4388), .A2(net_4387) );
HA_X1 inst_6709 ( .CO(net_1749), .S(net_1486), .A(net_1284), .B(net_838) );
INV_X4 inst_5805 ( .A(net_7589), .ZN(net_623) );
DFFS_X1 inst_6939 ( .D(net_6145), .CK(net_13649), .SN(x6501), .Q(x729) );
NAND2_X2 inst_4641 ( .ZN(net_2802), .A2(net_2418), .A1(net_2114) );
DFFR_X2 inst_7056 ( .QN(net_7499), .D(net_4820), .CK(net_16672), .RN(x6501) );
CLKBUF_X2 inst_11038 ( .A(net_9570), .Z(net_10886) );
SDFF_X2 inst_460 ( .SI(net_8464), .Q(net_8464), .SE(net_3983), .D(net_3974), .CK(net_12281) );
CLKBUF_X2 inst_10877 ( .A(net_10724), .Z(net_10725) );
SDFF_X2 inst_1455 ( .SI(net_7273), .Q(net_7050), .D(net_7050), .SE(net_6280), .CK(net_14137) );
DFFR_X2 inst_7135 ( .QN(net_6398), .D(net_2982), .CK(net_15693), .RN(x6501) );
SDFFR_X2 inst_2497 ( .SI(net_2539), .SE(net_2220), .Q(net_402), .D(net_402), .CK(net_14798), .RN(x6501) );
NAND4_X2 inst_3660 ( .A4(net_6012), .A1(net_6011), .ZN(net_4605), .A2(net_4132), .A3(net_4131) );
CLKBUF_X2 inst_16975 ( .A(net_15302), .Z(net_16823) );
CLKBUF_X2 inst_15678 ( .A(net_9278), .Z(net_15526) );
CLKBUF_X2 inst_16274 ( .A(net_16121), .Z(net_16122) );
NAND2_X2 inst_4230 ( .A1(net_7019), .A2(net_5249), .ZN(net_5230) );
CLKBUF_X2 inst_15316 ( .A(net_15163), .Z(net_15164) );
CLKBUF_X2 inst_16771 ( .A(net_16618), .Z(net_16619) );
INV_X4 inst_5571 ( .A(net_7363), .ZN(net_2123) );
CLKBUF_X2 inst_13455 ( .A(net_13302), .Z(net_13303) );
SDFF_X2 inst_950 ( .SI(net_7334), .Q(net_6708), .D(net_6708), .SE(net_3125), .CK(net_12051) );
NAND3_X2 inst_3955 ( .ZN(net_3148), .A1(net_3036), .A2(net_2097), .A3(net_1534) );
SDFF_X2 inst_1218 ( .Q(net_7942), .D(net_7942), .SE(net_2755), .SI(net_2721), .CK(net_15787) );
AOI22_X2 inst_8458 ( .B1(net_6671), .A1(net_6638), .A2(net_6213), .B2(net_6138), .ZN(net_3482) );
INV_X2 inst_6414 ( .ZN(net_1589), .A(net_862) );
CLKBUF_X2 inst_15842 ( .A(net_11523), .Z(net_15690) );
CLKBUF_X2 inst_9541 ( .A(net_9388), .Z(net_9389) );
XOR2_X1 inst_101 ( .A(net_1211), .Z(net_1207), .B(net_1206) );
CLKBUF_X2 inst_17696 ( .A(net_10832), .Z(net_17544) );
CLKBUF_X2 inst_14033 ( .A(net_13880), .Z(net_13881) );
NOR2_X2 inst_3555 ( .A2(net_8217), .ZN(net_2274), .A1(net_1317) );
CLKBUF_X2 inst_10234 ( .A(net_9357), .Z(net_10082) );
CLKBUF_X2 inst_14377 ( .A(net_13233), .Z(net_14225) );
CLKBUF_X2 inst_11388 ( .A(net_10461), .Z(net_11236) );
NAND2_X2 inst_4722 ( .A1(net_7372), .ZN(net_1970), .A2(net_1784) );
SDFF_X2 inst_510 ( .Q(net_8863), .D(net_8863), .SI(net_3962), .SE(net_3936), .CK(net_10174) );
CLKBUF_X2 inst_12194 ( .A(net_12041), .Z(net_12042) );
INV_X2 inst_6505 ( .A(net_7437), .ZN(net_537) );
SDFF_X2 inst_1677 ( .SI(net_7747), .Q(net_7747), .D(net_2573), .SE(net_2560), .CK(net_18037) );
SDFF_X2 inst_830 ( .SI(net_8491), .Q(net_8491), .D(net_3946), .SE(net_3884), .CK(net_10694) );
AOI22_X2 inst_8433 ( .B1(net_6731), .A1(net_6698), .B2(net_6202), .A2(net_3520), .ZN(net_3508) );
CLKBUF_X2 inst_15646 ( .A(net_15493), .Z(net_15494) );
OR2_X2 inst_2878 ( .ZN(net_3312), .A2(net_3311), .A1(net_3217) );
SDFFR_X2 inst_2494 ( .Q(net_8998), .D(net_8998), .SI(net_2602), .SE(net_2562), .CK(net_14532), .RN(x6501) );
SDFF_X2 inst_776 ( .SI(net_8334), .Q(net_8334), .D(net_3961), .SE(net_3880), .CK(net_10149) );
CLKBUF_X2 inst_18480 ( .A(net_18327), .Z(net_18328) );
SDFFR_X2 inst_2526 ( .D(net_7366), .SE(net_2387), .SI(net_281), .Q(net_281), .CK(net_13671), .RN(x6501) );
INV_X8 inst_5047 ( .A(net_6142), .ZN(net_6141) );
CLKBUF_X2 inst_10787 ( .A(net_10634), .Z(net_10635) );
INV_X4 inst_5313 ( .ZN(net_1473), .A(net_1104) );
SDFF_X2 inst_1972 ( .D(net_7272), .SI(net_7009), .Q(net_7009), .SE(net_6277), .CK(net_16796) );
SDFF_X2 inst_558 ( .Q(net_8672), .D(net_8672), .SI(net_3965), .SE(net_3935), .CK(net_12453) );
INV_X32 inst_6167 ( .ZN(net_5166), .A(net_4818) );
CLKBUF_X2 inst_12704 ( .A(net_12551), .Z(net_12552) );
CLKBUF_X2 inst_10591 ( .A(net_9781), .Z(net_10439) );
SDFF_X2 inst_389 ( .Q(net_8817), .D(net_8817), .SI(net_3980), .SE(net_3964), .CK(net_10741) );
INV_X4 inst_5179 ( .ZN(net_2996), .A(net_2911) );
CLKBUF_X2 inst_14301 ( .A(net_14148), .Z(net_14149) );
CLKBUF_X2 inst_13460 ( .A(net_13250), .Z(net_13308) );
SDFFR_X1 inst_2712 ( .QN(net_6818), .SE(net_6267), .SI(net_4617), .D(net_4373), .CK(net_11780), .RN(x6501) );
CLKBUF_X2 inst_16257 ( .A(net_11598), .Z(net_16105) );
CLKBUF_X2 inst_10252 ( .A(net_9381), .Z(net_10100) );
INV_X4 inst_6152 ( .ZN(net_6179), .A(net_2002) );
AOI222_X1 inst_8650 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3916), .B1(net_2151), .C1(net_2150), .A1(x13853) );
SDFF_X2 inst_1382 ( .SI(net_7295), .Q(net_7112), .D(net_7112), .SE(net_6278), .CK(net_18216) );
AOI221_X2 inst_8841 ( .B1(net_8049), .C1(net_7845), .B2(net_6107), .ZN(net_6027), .C2(net_4400), .A(net_4281) );
OR3_X4 inst_2795 ( .ZN(net_4409), .A1(net_4408), .A2(net_4407), .A3(net_4406) );
INV_X4 inst_5266 ( .A(net_2400), .ZN(net_2315) );
NAND2_X2 inst_4766 ( .ZN(net_1876), .A2(net_1681), .A1(net_716) );
NAND2_X2 inst_4445 ( .A1(net_6845), .A2(net_5016), .ZN(net_4982) );
INV_X4 inst_5895 ( .A(net_7607), .ZN(net_2230) );
CLKBUF_X2 inst_16545 ( .A(net_16392), .Z(net_16393) );
CLKBUF_X2 inst_17726 ( .A(net_17573), .Z(net_17574) );
CLKBUF_X2 inst_15898 ( .A(net_15745), .Z(net_15746) );
CLKBUF_X2 inst_11785 ( .A(net_11632), .Z(net_11633) );
CLKBUF_X2 inst_9977 ( .A(net_9818), .Z(net_9825) );
CLKBUF_X2 inst_12866 ( .A(net_12713), .Z(net_12714) );
CLKBUF_X2 inst_12766 ( .A(net_11219), .Z(net_12614) );
AOI22_X2 inst_8365 ( .B1(net_8592), .A1(net_8481), .A2(net_6263), .B2(net_6262), .ZN(net_3683) );
CLKBUF_X2 inst_14195 ( .A(net_11038), .Z(net_14043) );
CLKBUF_X2 inst_19108 ( .A(net_18955), .Z(net_18956) );
DFFR_X2 inst_7105 ( .QN(net_7344), .D(net_6196), .CK(net_9568), .RN(x6501) );
CLKBUF_X2 inst_10843 ( .A(net_10690), .Z(net_10691) );
CLKBUF_X2 inst_18064 ( .A(net_17911), .Z(net_17912) );
CLKBUF_X2 inst_16789 ( .A(net_13253), .Z(net_16637) );
CLKBUF_X2 inst_11613 ( .A(net_11460), .Z(net_11461) );
CLKBUF_X2 inst_11133 ( .A(net_10980), .Z(net_10981) );
CLKBUF_X2 inst_16067 ( .A(net_15914), .Z(net_15915) );
CLKBUF_X2 inst_11724 ( .A(net_10276), .Z(net_11572) );
CLKBUF_X2 inst_19015 ( .A(net_18862), .Z(net_18863) );
CLKBUF_X2 inst_17837 ( .A(net_14684), .Z(net_17685) );
CLKBUF_X2 inst_13321 ( .A(net_13168), .Z(net_13169) );
CLKBUF_X2 inst_9446 ( .A(net_9293), .Z(net_9294) );
CLKBUF_X2 inst_18685 ( .A(net_18532), .Z(net_18533) );
CLKBUF_X2 inst_13467 ( .A(net_13314), .Z(net_13315) );
NAND2_X2 inst_4212 ( .A1(net_7010), .ZN(net_5250), .A2(net_5249) );
CLKBUF_X2 inst_15257 ( .A(net_15104), .Z(net_15105) );
CLKBUF_X2 inst_15716 ( .A(net_15563), .Z(net_15564) );
CLKBUF_X2 inst_11231 ( .A(net_11078), .Z(net_11079) );
CLKBUF_X2 inst_12912 ( .A(net_12759), .Z(net_12760) );
CLKBUF_X2 inst_11759 ( .A(net_11606), .Z(net_11607) );
CLKBUF_X2 inst_9594 ( .A(net_9441), .Z(net_9442) );
CLKBUF_X2 inst_16238 ( .A(net_9577), .Z(net_16086) );
SDFFR_X2 inst_2309 ( .SE(net_2260), .Q(net_363), .D(net_363), .CK(net_11476), .RN(x6501), .SI(x1855) );
CLKBUF_X2 inst_15011 ( .A(net_10332), .Z(net_14859) );
CLKBUF_X2 inst_16285 ( .A(net_16132), .Z(net_16133) );
DFFR_X2 inst_7196 ( .QN(net_8954), .D(net_2419), .CK(net_15193), .RN(x6501) );
CLKBUF_X2 inst_18225 ( .A(net_18072), .Z(net_18073) );
CLKBUF_X2 inst_11283 ( .A(net_11130), .Z(net_11131) );
SDFFR_X2 inst_2603 ( .D(net_7368), .Q(net_7265), .SI(net_1854), .SE(net_1327), .CK(net_14679), .RN(x6501) );
CLKBUF_X2 inst_15792 ( .A(net_15639), .Z(net_15640) );
CLKBUF_X2 inst_11335 ( .A(net_11182), .Z(net_11183) );
NAND2_X2 inst_4603 ( .A2(net_6127), .ZN(net_2850), .A1(net_2532) );
CLKBUF_X2 inst_9339 ( .A(net_9186), .Z(net_9187) );
SDFFR_X2 inst_2153 ( .Q(net_8279), .D(net_3241), .SE(net_2996), .SI(net_1212), .CK(net_18442), .RN(x6501) );
CLKBUF_X2 inst_18808 ( .A(net_18655), .Z(net_18656) );
CLKBUF_X2 inst_11271 ( .A(net_11118), .Z(net_11119) );
CLKBUF_X2 inst_11904 ( .A(net_11751), .Z(net_11752) );
CLKBUF_X2 inst_11798 ( .A(net_11645), .Z(net_11646) );
CLKBUF_X2 inst_18759 ( .A(net_18606), .Z(net_18607) );
CLKBUF_X2 inst_16996 ( .A(net_16843), .Z(net_16844) );
INV_X4 inst_5494 ( .ZN(net_856), .A(net_718) );
CLKBUF_X2 inst_10586 ( .A(net_10433), .Z(net_10434) );
INV_X4 inst_5441 ( .ZN(net_1140), .A(net_821) );
CLKBUF_X2 inst_9906 ( .A(net_9753), .Z(net_9754) );
DFFS_X2 inst_6874 ( .QN(net_7651), .D(net_3900), .CK(net_12667), .SN(x6501) );
NOR2_X2 inst_3485 ( .ZN(net_2124), .A1(net_2123), .A2(net_2122) );
INV_X4 inst_5854 ( .A(net_7441), .ZN(net_1037) );
AOI222_X2 inst_8587 ( .B2(net_6782), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5817), .A1(net_4208), .C1(x2451) );
AOI222_X1 inst_8680 ( .A2(net_3296), .B2(net_3295), .C2(net_3294), .ZN(net_3293), .A1(net_3292), .C1(net_3032), .B1(net_1465) );
HA_X1 inst_6678 ( .S(net_3102), .CO(net_3101), .B(net_3046), .A(x2594) );
CLKBUF_X2 inst_17646 ( .A(net_12639), .Z(net_17494) );
CLKBUF_X2 inst_16451 ( .A(net_16298), .Z(net_16299) );
CLKBUF_X2 inst_9616 ( .A(net_9463), .Z(net_9464) );
CLKBUF_X2 inst_12798 ( .A(net_12617), .Z(net_12646) );
CLKBUF_X2 inst_16367 ( .A(net_16214), .Z(net_16215) );
DFFR_X2 inst_7011 ( .QN(net_6294), .D(net_5761), .CK(net_16746), .RN(x6501) );
DFFR_X2 inst_7201 ( .D(net_2366), .QN(net_226), .CK(net_17798), .RN(x6501) );
CLKBUF_X2 inst_11049 ( .A(net_10896), .Z(net_10897) );
CLKBUF_X2 inst_9649 ( .A(net_9470), .Z(net_9497) );
CLKBUF_X2 inst_9320 ( .A(net_9167), .Z(net_9168) );
SDFF_X2 inst_620 ( .SI(net_8531), .Q(net_8531), .SE(net_3979), .D(net_3945), .CK(net_11088) );
INV_X2 inst_6496 ( .A(net_7624), .ZN(net_549) );
OAI21_X2 inst_3118 ( .A(net_5955), .ZN(net_2331), .B2(net_1642), .B1(net_1205) );
INV_X2 inst_6401 ( .ZN(net_1604), .A(net_1152) );
CLKBUF_X2 inst_18944 ( .A(net_18353), .Z(net_18792) );
DFFS_X2 inst_6869 ( .QN(net_6808), .D(net_4620), .CK(net_11804), .SN(x6501) );
CLKBUF_X2 inst_14597 ( .A(net_14444), .Z(net_14445) );
CLKBUF_X2 inst_14514 ( .A(net_14361), .Z(net_14362) );
SDFF_X2 inst_1409 ( .SI(net_7276), .Q(net_7053), .D(net_7053), .SE(net_6280), .CK(net_17389) );
CLKBUF_X2 inst_10757 ( .A(net_9951), .Z(net_10605) );
CLKBUF_X2 inst_11570 ( .A(net_11417), .Z(net_11418) );
CLKBUF_X2 inst_13752 ( .A(net_13599), .Z(net_13600) );
CLKBUF_X2 inst_15613 ( .A(net_9679), .Z(net_15461) );
CLKBUF_X2 inst_13509 ( .A(net_13356), .Z(net_13357) );
OAI21_X2 inst_2996 ( .B2(net_5902), .ZN(net_5897), .A(net_5819), .B1(net_671) );
INV_X8 inst_5037 ( .ZN(net_6094), .A(net_1682) );
CLKBUF_X2 inst_10601 ( .A(net_9145), .Z(net_10449) );
CLKBUF_X2 inst_16261 ( .A(net_16108), .Z(net_16109) );
CLKBUF_X2 inst_16762 ( .A(net_16609), .Z(net_16610) );
CLKBUF_X2 inst_11946 ( .A(net_11181), .Z(net_11794) );
CLKBUF_X2 inst_9517 ( .A(net_9364), .Z(net_9365) );
CLKBUF_X2 inst_14002 ( .A(net_13828), .Z(net_13850) );
AOI221_X2 inst_8763 ( .C2(net_6130), .B2(net_5535), .ZN(net_5469), .A(net_4945), .C1(net_1389), .B1(net_464) );
XOR2_X2 inst_4 ( .Z(net_3116), .A(net_2978), .B(x2746) );
NAND4_X2 inst_3795 ( .ZN(net_3631), .A1(net_3508), .A2(net_3507), .A3(net_3506), .A4(net_3505) );
CLKBUF_X2 inst_18323 ( .A(net_18170), .Z(net_18171) );
NOR3_X2 inst_3272 ( .A1(net_2415), .ZN(net_2414), .A3(net_2397), .A2(net_1864) );
CLKBUF_X2 inst_9846 ( .A(net_9693), .Z(net_9694) );
CLKBUF_X2 inst_9455 ( .A(net_9302), .Z(net_9303) );
CLKBUF_X2 inst_10494 ( .A(net_10341), .Z(net_10342) );
CLKBUF_X2 inst_14232 ( .A(net_14079), .Z(net_14080) );
SDFF_X2 inst_1866 ( .D(net_7266), .SI(net_6923), .Q(net_6923), .SE(net_6281), .CK(net_14343) );
CLKBUF_X2 inst_15230 ( .A(net_11179), .Z(net_15078) );
AOI221_X2 inst_8795 ( .C2(net_6187), .B2(net_5609), .ZN(net_4900), .A(net_4898), .B1(net_372), .C1(net_196) );
SDFF_X2 inst_1878 ( .D(net_7286), .SI(net_6983), .Q(net_6983), .SE(net_6283), .CK(net_17669) );
INV_X4 inst_5136 ( .A(net_3552), .ZN(net_3549) );
CLKBUF_X2 inst_18240 ( .A(net_18087), .Z(net_18088) );
INV_X4 inst_6016 ( .A(net_7392), .ZN(net_1650) );
CLKBUF_X2 inst_16459 ( .A(net_16306), .Z(net_16307) );
CLKBUF_X2 inst_10290 ( .A(net_10137), .Z(net_10138) );
SDFF_X2 inst_765 ( .Q(net_8780), .D(net_8780), .SI(net_3980), .SE(net_3879), .CK(net_13331) );
CLKBUF_X2 inst_10790 ( .A(net_9607), .Z(net_10638) );
CLKBUF_X2 inst_9870 ( .A(net_9717), .Z(net_9718) );
CLKBUF_X2 inst_17434 ( .A(net_16250), .Z(net_17282) );
CLKBUF_X2 inst_10664 ( .A(net_9875), .Z(net_10512) );
CLKBUF_X2 inst_14247 ( .A(net_14094), .Z(net_14095) );
NOR2_X2 inst_3422 ( .ZN(net_3296), .A2(net_3294), .A1(net_3068) );
CLKBUF_X2 inst_13266 ( .A(net_10794), .Z(net_13114) );
NAND4_X2 inst_3832 ( .ZN(net_2295), .A2(net_2024), .A1(net_2023), .A4(net_1416), .A3(net_1386) );
INV_X2 inst_6618 ( .ZN(net_6212), .A(net_6209) );
NAND2_X4 inst_4039 ( .A1(net_6258), .ZN(net_6128), .A2(net_5990) );
OAI221_X2 inst_2967 ( .C1(net_8945), .ZN(net_2651), .B2(net_2650), .C2(net_2649), .A(net_2478), .B1(net_1488) );
CLKBUF_X2 inst_16681 ( .A(net_16528), .Z(net_16529) );
CLKBUF_X2 inst_13279 ( .A(net_10950), .Z(net_13127) );
INV_X4 inst_5674 ( .A(net_8890), .ZN(net_1156) );
AND4_X4 inst_9029 ( .ZN(net_1904), .A2(net_1723), .A3(net_1722), .A4(net_1373), .A1(net_632) );
CLKBUF_X2 inst_14873 ( .A(net_14720), .Z(net_14721) );
SDFF_X2 inst_699 ( .Q(net_8437), .D(net_8437), .SI(net_3952), .SE(net_3934), .CK(net_10348) );
AOI22_X2 inst_8377 ( .B1(net_8745), .A1(net_8375), .A2(net_3867), .B2(net_3866), .ZN(net_3671) );
CLKBUF_X2 inst_9921 ( .A(net_9768), .Z(net_9769) );
CLKBUF_X2 inst_18025 ( .A(net_17872), .Z(net_17873) );
CLKBUF_X2 inst_9514 ( .A(net_9076), .Z(net_9362) );
CLKBUF_X2 inst_13823 ( .A(net_13670), .Z(net_13671) );
CLKBUF_X2 inst_18644 ( .A(net_17735), .Z(net_18492) );
CLKBUF_X2 inst_14880 ( .A(net_14727), .Z(net_14728) );
CLKBUF_X2 inst_13144 ( .A(net_12991), .Z(net_12992) );
SDFFR_X2 inst_2426 ( .SE(net_2678), .D(net_2675), .SI(net_448), .Q(net_448), .CK(net_13845), .RN(x6501) );
CLKBUF_X2 inst_14211 ( .A(net_14058), .Z(net_14059) );
INV_X2 inst_6377 ( .A(net_1372), .ZN(net_1354) );
CLKBUF_X2 inst_14528 ( .A(net_10752), .Z(net_14376) );
CLKBUF_X2 inst_18304 ( .A(net_18151), .Z(net_18152) );
CLKBUF_X2 inst_18260 ( .A(net_14961), .Z(net_18108) );
CLKBUF_X2 inst_17547 ( .A(net_17394), .Z(net_17395) );
SDFF_X2 inst_1485 ( .SI(net_7296), .Q(net_7073), .D(net_7073), .SE(net_6280), .CK(net_15453) );
CLKBUF_X2 inst_17283 ( .A(net_9900), .Z(net_17131) );
CLKBUF_X2 inst_12259 ( .A(net_12106), .Z(net_12107) );
SDFF_X2 inst_750 ( .Q(net_8789), .D(net_8789), .SI(net_3962), .SE(net_3879), .CK(net_12955) );
XNOR2_X2 inst_317 ( .ZN(net_947), .B(net_943), .A(net_206) );
CLKBUF_X2 inst_10561 ( .A(net_10408), .Z(net_10409) );
AOI21_X2 inst_8947 ( .A(net_5783), .ZN(net_5677), .B1(net_5473), .B2(net_5269) );
XNOR2_X2 inst_278 ( .A(net_6833), .ZN(net_1030), .B(net_1029) );
NAND2_X2 inst_4429 ( .A1(net_6867), .A2(net_5016), .ZN(net_4998) );
SDFF_X2 inst_467 ( .SI(net_8472), .Q(net_8472), .SE(net_3983), .D(net_3941), .CK(net_12905) );
CLKBUF_X2 inst_16117 ( .A(net_15964), .Z(net_15965) );
NAND4_X2 inst_3677 ( .A4(net_6026), .A1(net_6025), .ZN(net_4588), .A2(net_4029), .A3(net_4028) );
NOR2_X2 inst_3456 ( .ZN(net_2971), .A2(net_2691), .A1(net_1442) );
CLKBUF_X2 inst_17370 ( .A(net_17217), .Z(net_17218) );
OAI221_X2 inst_2963 ( .C1(net_7353), .ZN(net_3066), .C2(net_3064), .B2(net_3063), .A(net_2883), .B1(net_2213) );
AOI22_X2 inst_7923 ( .A1(net_8992), .A2(net_5456), .B2(net_5260), .ZN(net_4458), .B1(net_4457) );
CLKBUF_X2 inst_10535 ( .A(net_10382), .Z(net_10383) );
SDFF_X2 inst_1329 ( .SI(net_7671), .Q(net_7671), .SE(net_2714), .D(net_2585), .CK(net_18565) );
SDFF_X2 inst_1204 ( .Q(net_7944), .D(net_7944), .SE(net_2755), .SI(net_2705), .CK(net_18594) );
AOI222_X1 inst_8687 ( .A1(net_6459), .A2(net_3296), .B2(net_3295), .C2(net_3294), .ZN(net_3283), .C1(net_3282), .B1(net_2876) );
NAND2_X2 inst_4066 ( .ZN(net_5873), .A2(net_5767), .A1(net_3584) );
CLKBUF_X2 inst_17974 ( .A(net_17821), .Z(net_17822) );
CLKBUF_X2 inst_13568 ( .A(net_11823), .Z(net_13416) );
CLKBUF_X2 inst_13158 ( .A(net_13005), .Z(net_13006) );
CLKBUF_X2 inst_10162 ( .A(net_10009), .Z(net_10010) );
CLKBUF_X2 inst_17687 ( .A(net_9964), .Z(net_17535) );
CLKBUF_X2 inst_11015 ( .A(net_10862), .Z(net_10863) );
CLKBUF_X2 inst_11718 ( .A(net_11565), .Z(net_11566) );
SDFFR_X2 inst_2618 ( .Q(net_7374), .D(net_7374), .SE(net_1136), .CK(net_18628), .RN(x6501), .SI(x4788) );
CLKBUF_X2 inst_15065 ( .A(net_14912), .Z(net_14913) );
CLKBUF_X2 inst_10952 ( .A(net_10799), .Z(net_10800) );
MUX2_X2 inst_4950 ( .A(net_7374), .S(net_2376), .Z(net_2374), .B(net_888) );
CLKBUF_X2 inst_14726 ( .A(net_14573), .Z(net_14574) );
AOI221_X2 inst_8853 ( .B1(net_8878), .C1(net_8323), .B2(net_6252), .ZN(net_6227), .C2(net_4345), .A(net_4249) );
CLKBUF_X2 inst_11443 ( .A(net_9565), .Z(net_11291) );
CLKBUF_X2 inst_9241 ( .A(net_9088), .Z(net_9089) );
CLKBUF_X2 inst_19053 ( .A(net_18900), .Z(net_18901) );
CLKBUF_X2 inst_17943 ( .A(net_17790), .Z(net_17791) );
CLKBUF_X2 inst_16916 ( .A(net_10842), .Z(net_16764) );
CLKBUF_X2 inst_14428 ( .A(net_14275), .Z(net_14276) );
SDFF_X2 inst_1729 ( .Q(net_7976), .D(net_7976), .SI(net_2721), .SE(net_2542), .CK(net_15820) );
AOI22_X2 inst_8346 ( .B1(net_8885), .A1(net_8330), .B2(net_6252), .A2(net_4345), .ZN(net_3701) );
CLKBUF_X2 inst_13175 ( .A(net_13022), .Z(net_13023) );
INV_X4 inst_6126 ( .A(net_8259), .ZN(net_2989) );
DFFR_X2 inst_6996 ( .QN(net_6297), .D(net_5842), .CK(net_16755), .RN(x6501) );
CLKBUF_X2 inst_13576 ( .A(net_9841), .Z(net_13424) );
CLKBUF_X2 inst_15202 ( .A(net_15049), .Z(net_15050) );
NAND2_X2 inst_4648 ( .A1(net_2346), .A2(net_2341), .ZN(net_2340) );
CLKBUF_X2 inst_10469 ( .A(net_9422), .Z(net_10317) );
CLKBUF_X2 inst_10297 ( .A(net_9616), .Z(net_10145) );
CLKBUF_X2 inst_11460 ( .A(net_11307), .Z(net_11308) );
XNOR2_X2 inst_165 ( .ZN(net_1828), .A(net_1603), .B(net_1495) );
NAND4_X2 inst_3733 ( .ZN(net_4297), .A1(net_4118), .A2(net_4117), .A3(net_4116), .A4(net_4115) );
INV_X4 inst_5376 ( .ZN(net_1378), .A(net_1342) );
SDFF_X2 inst_1176 ( .SI(net_7319), .Q(net_6594), .D(net_6594), .SE(net_3069), .CK(net_9832) );
CLKBUF_X2 inst_17102 ( .A(net_16949), .Z(net_16950) );
CLKBUF_X2 inst_12537 ( .A(net_9739), .Z(net_12385) );
AOI22_X2 inst_8159 ( .A1(net_7951), .B1(net_7781), .A2(net_6092), .B2(net_6091), .ZN(net_3993) );
CLKBUF_X2 inst_18127 ( .A(net_17974), .Z(net_17975) );
CLKBUF_X2 inst_12696 ( .A(net_12458), .Z(net_12544) );
INV_X4 inst_5450 ( .A(net_1063), .ZN(net_806) );
CLKBUF_X2 inst_15706 ( .A(net_15553), .Z(net_15554) );
CLKBUF_X2 inst_11340 ( .A(net_10071), .Z(net_11188) );
NAND2_X2 inst_4172 ( .ZN(net_5337), .A1(net_5195), .A2(net_4990) );
CLKBUF_X2 inst_13388 ( .A(net_13235), .Z(net_13236) );
SDFFR_X2 inst_2605 ( .D(net_7372), .Q(net_7269), .SI(net_1809), .SE(net_1327), .CK(net_17513), .RN(x6501) );
CLKBUF_X2 inst_14423 ( .A(net_14219), .Z(net_14271) );
CLKBUF_X2 inst_14147 ( .A(net_11610), .Z(net_13995) );
CLKBUF_X2 inst_13759 ( .A(net_11005), .Z(net_13607) );
DFFR_X2 inst_7252 ( .QN(net_7304), .D(net_2044), .CK(net_15043), .RN(x6501) );
CLKBUF_X2 inst_13717 ( .A(net_13564), .Z(net_13565) );
SDFFR_X1 inst_2703 ( .SI(net_7535), .SE(net_5043), .CK(net_11928), .RN(x6501), .Q(x4115), .D(x4115) );
CLKBUF_X2 inst_17464 ( .A(net_17311), .Z(net_17312) );
CLKBUF_X2 inst_13857 ( .A(net_13704), .Z(net_13705) );
CLKBUF_X2 inst_9784 ( .A(net_9631), .Z(net_9632) );
XNOR2_X2 inst_143 ( .ZN(net_2302), .B(net_2230), .A(net_2229) );
CLKBUF_X2 inst_15958 ( .A(net_11065), .Z(net_15806) );
CLKBUF_X2 inst_16698 ( .A(net_16545), .Z(net_16546) );
INV_X4 inst_5286 ( .ZN(net_1984), .A(net_1379) );
INV_X2 inst_6260 ( .ZN(net_4637), .A(net_4527) );
NAND2_X2 inst_4272 ( .A1(net_7038), .A2(net_5249), .ZN(net_5188) );
CLKBUF_X2 inst_16403 ( .A(net_16250), .Z(net_16251) );
CLKBUF_X2 inst_16878 ( .A(net_12778), .Z(net_16726) );
SDFFR_X2 inst_2337 ( .SE(net_2260), .Q(net_369), .D(net_369), .CK(net_11459), .RN(x6501), .SI(x1690) );
NOR4_X2 inst_3250 ( .A3(net_5971), .A4(net_5970), .A1(net_5969), .A2(net_5968), .ZN(net_2393) );
CLKBUF_X2 inst_15052 ( .A(net_14899), .Z(net_14900) );
CLKBUF_X2 inst_9357 ( .A(net_9105), .Z(net_9205) );
SDFF_X2 inst_1778 ( .SI(net_8072), .Q(net_8072), .D(net_2715), .SE(net_2508), .CK(net_14246) );
CLKBUF_X2 inst_18991 ( .A(net_18838), .Z(net_18839) );
CLKBUF_X2 inst_16158 ( .A(net_11942), .Z(net_16006) );
CLKBUF_X2 inst_12132 ( .A(net_11979), .Z(net_11980) );
AOI22_X2 inst_8091 ( .A1(net_7972), .B1(net_7802), .A2(net_6092), .B2(net_6091), .ZN(net_4055) );
SDFF_X2 inst_1736 ( .Q(net_8130), .D(net_8130), .SI(net_2590), .SE(net_2541), .CK(net_15572) );
SDFF_X2 inst_1040 ( .SI(net_7339), .Q(net_6713), .D(net_6713), .SE(net_3125), .CK(net_11896) );
NAND2_X4 inst_4027 ( .A2(net_6178), .A1(net_5989), .ZN(net_3081) );
CLKBUF_X2 inst_16648 ( .A(net_16495), .Z(net_16496) );
CLKBUF_X2 inst_15218 ( .A(net_15065), .Z(net_15066) );
AND2_X2 inst_9158 ( .ZN(net_2830), .A1(net_2829), .A2(net_2828) );
INV_X4 inst_6009 ( .A(net_8946), .ZN(net_662) );
INV_X8 inst_5042 ( .ZN(net_6102), .A(net_3556) );
CLKBUF_X2 inst_17032 ( .A(net_12281), .Z(net_16880) );
CLKBUF_X2 inst_16218 ( .A(net_16065), .Z(net_16066) );
OAI21_X2 inst_3146 ( .B2(net_2048), .ZN(net_2026), .A(net_2025), .B1(net_1125) );
CLKBUF_X2 inst_10246 ( .A(net_9462), .Z(net_10094) );
DFFR_X2 inst_7303 ( .QN(net_8269), .D(net_8265), .CK(net_18491), .RN(x6501) );
CLKBUF_X2 inst_11651 ( .A(net_11498), .Z(net_11499) );
SDFF_X2 inst_2056 ( .SI(net_7797), .Q(net_7797), .D(net_2711), .SE(net_2459), .CK(net_14233) );
SDFFR_X2 inst_2116 ( .SI(net_7179), .Q(net_7179), .D(net_6430), .SE(net_4362), .CK(net_13579), .RN(x6501) );
OR2_X4 inst_2825 ( .A2(net_6158), .ZN(net_4490), .A1(net_3927) );
INV_X4 inst_5071 ( .ZN(net_5857), .A(net_5811) );
CLKBUF_X2 inst_17135 ( .A(net_16982), .Z(net_16983) );
NAND2_X4 inst_4031 ( .ZN(net_3071), .A1(net_2905), .A2(net_2903) );
CLKBUF_X2 inst_16607 ( .A(net_16454), .Z(net_16455) );
CLKBUF_X2 inst_15370 ( .A(net_12660), .Z(net_15218) );
AOI22_X2 inst_8135 ( .A1(net_7948), .B1(net_7778), .A2(net_6092), .B2(net_6091), .ZN(net_4015) );
SDFF_X2 inst_346 ( .SI(net_8474), .Q(net_8474), .SE(net_3983), .D(net_3952), .CK(net_12912) );
AOI221_X2 inst_8755 ( .C1(net_7512), .ZN(net_5536), .B2(net_5535), .C2(net_5260), .A(net_5021), .B1(net_471) );
CLKBUF_X2 inst_10711 ( .A(net_10558), .Z(net_10559) );
CLKBUF_X2 inst_12058 ( .A(net_11905), .Z(net_11906) );
INV_X2 inst_6195 ( .A(net_6790), .ZN(net_5731) );
CLKBUF_X2 inst_9777 ( .A(net_9624), .Z(net_9625) );
CLKBUF_X2 inst_11347 ( .A(net_10296), .Z(net_11195) );
CLKBUF_X2 inst_12972 ( .A(net_12819), .Z(net_12820) );
NAND3_X2 inst_3929 ( .ZN(net_5586), .A1(net_5460), .A3(net_4768), .A2(net_4573) );
AOI221_X2 inst_8856 ( .B1(net_8886), .C1(net_8331), .B2(net_6252), .ZN(net_6237), .C2(net_4345), .A(net_4240) );
CLKBUF_X2 inst_12312 ( .A(net_9683), .Z(net_12160) );
CLKBUF_X2 inst_10506 ( .A(net_10353), .Z(net_10354) );
NAND4_X2 inst_3852 ( .ZN(net_1560), .A3(net_1025), .A2(net_1006), .A4(net_986), .A1(net_953) );
CLKBUF_X2 inst_18549 ( .A(net_18396), .Z(net_18397) );
CLKBUF_X2 inst_15131 ( .A(net_14978), .Z(net_14979) );
CLKBUF_X2 inst_14168 ( .A(net_14015), .Z(net_14016) );
SDFF_X2 inst_1051 ( .SI(net_7336), .Q(net_6677), .D(net_6677), .SE(net_3126), .CK(net_9481) );
SDFFR_X2 inst_2566 ( .QN(net_6354), .SE(net_2147), .D(net_2126), .SI(net_1809), .CK(net_17526), .RN(x6501) );
CLKBUF_X2 inst_19024 ( .A(net_18871), .Z(net_18872) );
INV_X4 inst_6102 ( .A(net_7373), .ZN(net_1225) );
CLKBUF_X2 inst_18690 ( .A(net_11297), .Z(net_18538) );
CLKBUF_X2 inst_12901 ( .A(net_12748), .Z(net_12749) );
NOR2_X2 inst_3603 ( .A1(net_7519), .ZN(net_1526), .A2(net_740) );
CLKBUF_X2 inst_11076 ( .A(net_10923), .Z(net_10924) );
OAI21_X2 inst_3043 ( .B2(net_8240), .B1(net_4928), .ZN(net_4786), .A(net_3204) );
AOI22_X2 inst_8063 ( .A1(net_7969), .B1(net_7799), .A2(net_6092), .B2(net_6091), .ZN(net_4079) );
CLKBUF_X2 inst_13665 ( .A(net_13512), .Z(net_13513) );
INV_X4 inst_5752 ( .A(net_5972), .ZN(x3372) );
CLKBUF_X2 inst_14969 ( .A(net_14816), .Z(net_14817) );
CLKBUF_X2 inst_10548 ( .A(net_10302), .Z(net_10396) );
CLKBUF_X2 inst_13781 ( .A(net_13628), .Z(net_13629) );
CLKBUF_X2 inst_11360 ( .A(net_10494), .Z(net_11208) );
SDFF_X2 inst_573 ( .Q(net_8838), .D(net_8838), .SE(net_3964), .SI(net_3942), .CK(net_12627) );
AOI22_X4 inst_7736 ( .B2(net_8761), .A1(net_8391), .A2(net_3867), .B1(net_3866), .ZN(net_3789) );
CLKBUF_X2 inst_17735 ( .A(net_17582), .Z(net_17583) );
CLKBUF_X2 inst_17123 ( .A(net_9200), .Z(net_16971) );
CLKBUF_X2 inst_17757 ( .A(net_17604), .Z(net_17605) );
AND3_X4 inst_9041 ( .A3(net_6136), .ZN(net_2868), .A2(net_2540), .A1(net_1436) );
AOI22_X2 inst_8088 ( .B1(net_8074), .A1(net_7870), .B2(net_6107), .A2(net_4400), .ZN(net_4058) );
INV_X4 inst_5364 ( .A(net_2093), .ZN(net_1139) );
CLKBUF_X2 inst_18669 ( .A(net_18516), .Z(net_18517) );
NAND2_X2 inst_4245 ( .A1(net_6905), .A2(net_5247), .ZN(net_5215) );
CLKBUF_X2 inst_18169 ( .A(net_18016), .Z(net_18017) );
CLKBUF_X2 inst_17868 ( .A(net_17715), .Z(net_17716) );
CLKBUF_X2 inst_12391 ( .A(net_12238), .Z(net_12239) );
AOI21_X2 inst_8978 ( .B2(net_2146), .ZN(net_2105), .B1(net_2104), .A(net_2099) );
NOR2_X2 inst_3544 ( .A2(net_7417), .ZN(net_1678), .A1(net_1318) );
CLKBUF_X2 inst_10973 ( .A(net_10820), .Z(net_10821) );
CLKBUF_X2 inst_18871 ( .A(net_18718), .Z(net_18719) );
CLKBUF_X2 inst_17558 ( .A(net_9375), .Z(net_17406) );
AOI22_X2 inst_7970 ( .B1(net_8127), .A1(net_7889), .A2(net_6098), .B2(net_4190), .ZN(net_4159) );
CLKBUF_X2 inst_13607 ( .A(net_13454), .Z(net_13455) );
CLKBUF_X2 inst_17404 ( .A(net_17251), .Z(net_17252) );
CLKBUF_X2 inst_9362 ( .A(net_9107), .Z(net_9210) );
CLKBUF_X2 inst_18351 ( .A(net_18198), .Z(net_18199) );
INV_X2 inst_6367 ( .A(net_4394), .ZN(net_1729) );
CLKBUF_X2 inst_18656 ( .A(net_13373), .Z(net_18504) );
CLKBUF_X2 inst_15876 ( .A(net_15723), .Z(net_15724) );
INV_X4 inst_5553 ( .A(net_1252), .ZN(net_636) );
CLKBUF_X2 inst_11518 ( .A(net_11365), .Z(net_11366) );
INV_X4 inst_6111 ( .A(net_7166), .ZN(net_2031) );
NOR2_X2 inst_3522 ( .ZN(net_1888), .A1(net_1661), .A2(net_1621) );
CLKBUF_X2 inst_15795 ( .A(net_15642), .Z(net_15643) );
INV_X2 inst_6306 ( .ZN(net_3898), .A(net_3596) );
CLKBUF_X2 inst_14119 ( .A(net_13966), .Z(net_13967) );
CLKBUF_X2 inst_18475 ( .A(net_18322), .Z(net_18323) );
SDFF_X2 inst_1758 ( .Q(net_8127), .D(net_8127), .SI(net_2576), .SE(net_2541), .CK(net_16024) );
SDFF_X2 inst_1142 ( .SI(net_7321), .Q(net_6596), .D(net_6596), .SE(net_3069), .CK(net_12077) );
INV_X2 inst_6280 ( .ZN(net_4228), .A(net_3985) );
NAND4_X2 inst_3816 ( .ZN(net_3610), .A1(net_3423), .A2(net_3422), .A3(net_3421), .A4(net_3420) );
CLKBUF_X2 inst_11138 ( .A(net_10473), .Z(net_10986) );
CLKBUF_X2 inst_14914 ( .A(net_14761), .Z(net_14762) );
CLKBUF_X2 inst_15979 ( .A(net_15606), .Z(net_15827) );
CLKBUF_X2 inst_14772 ( .A(net_14619), .Z(net_14620) );
INV_X4 inst_5418 ( .ZN(net_1131), .A(net_860) );
CLKBUF_X2 inst_19152 ( .A(net_9577), .Z(net_19000) );
SDFF_X2 inst_1381 ( .SI(net_7734), .Q(net_7734), .D(net_2704), .SE(net_2559), .CK(net_14423) );
CLKBUF_X2 inst_15527 ( .A(net_13146), .Z(net_15375) );
SDFF_X2 inst_643 ( .SI(net_8525), .Q(net_8525), .SE(net_3979), .D(net_3947), .CK(net_12969) );
CLKBUF_X2 inst_12471 ( .A(net_12318), .Z(net_12319) );
CLKBUF_X2 inst_13726 ( .A(net_13573), .Z(net_13574) );
CLKBUF_X2 inst_9430 ( .A(net_9277), .Z(net_9278) );
CLKBUF_X2 inst_10745 ( .A(net_10592), .Z(net_10593) );
AOI22_X2 inst_7763 ( .B1(net_6990), .A1(net_6950), .A2(net_5443), .B2(net_5442), .ZN(net_5354) );
CLKBUF_X2 inst_12117 ( .A(net_11964), .Z(net_11965) );
CLKBUF_X2 inst_12220 ( .A(net_12067), .Z(net_12068) );
MUX2_X2 inst_4961 ( .A(net_7383), .S(net_2370), .Z(net_2362), .B(net_804) );
AOI222_X2 inst_8588 ( .B1(net_6187), .A2(net_6134), .C2(net_5538), .ZN(net_4921), .A1(net_1415), .C1(net_429), .B2(net_203) );
INV_X2 inst_6466 ( .A(net_7632), .ZN(net_577) );
CLKBUF_X2 inst_12165 ( .A(net_12012), .Z(net_12013) );
AOI22_X2 inst_8581 ( .ZN(net_1797), .A2(net_1344), .B2(net_757), .B1(net_689), .A1(x4869) );
INV_X4 inst_5447 ( .A(net_1253), .ZN(net_1080) );
INV_X2 inst_6371 ( .ZN(net_1820), .A(net_1659) );
CLKBUF_X2 inst_17538 ( .A(net_14340), .Z(net_17386) );
NAND2_X2 inst_4146 ( .ZN(net_5372), .A1(net_5110), .A2(net_5109) );
CLKBUF_X2 inst_12526 ( .A(net_12373), .Z(net_12374) );
CLKBUF_X2 inst_17220 ( .A(net_10253), .Z(net_17068) );
CLKBUF_X2 inst_12959 ( .A(net_12806), .Z(net_12807) );
SDFF_X2 inst_1997 ( .SI(net_7925), .Q(net_7925), .D(net_2719), .SE(net_2461), .CK(net_15568) );
DFFR_X2 inst_6971 ( .QN(net_7345), .D(net_5925), .CK(net_9583), .RN(x6501) );
CLKBUF_X2 inst_12669 ( .A(net_12516), .Z(net_12517) );
SDFFR_X2 inst_2297 ( .QN(net_7476), .SE(net_3354), .SI(net_3113), .CK(net_12160), .D(x13374), .RN(x6501) );
NAND4_X2 inst_3736 ( .ZN(net_4294), .A1(net_4100), .A2(net_4099), .A3(net_4098), .A4(net_4097) );
NOR2_X4 inst_3341 ( .A2(net_7415), .A1(net_7414), .ZN(net_1078) );
AOI22_X2 inst_8500 ( .B1(net_6548), .A1(net_6515), .A2(net_6137), .B2(net_6104), .ZN(net_3440) );
CLKBUF_X2 inst_13411 ( .A(net_13258), .Z(net_13259) );
INV_X2 inst_6374 ( .A(net_2912), .ZN(net_2906) );
CLKBUF_X2 inst_15296 ( .A(net_15143), .Z(net_15144) );
CLKBUF_X2 inst_14913 ( .A(net_14760), .Z(net_14761) );
SDFFR_X2 inst_2508 ( .Q(net_9000), .D(net_9000), .SI(net_4540), .SE(net_2562), .CK(net_14692), .RN(x6501) );
CLKBUF_X2 inst_10207 ( .A(net_9394), .Z(net_10055) );
CLKBUF_X2 inst_14642 ( .A(net_14489), .Z(net_14490) );
SDFF_X2 inst_773 ( .Q(net_8784), .D(net_8784), .SI(net_3947), .SE(net_3879), .CK(net_12954) );
CLKBUF_X2 inst_10776 ( .A(net_10623), .Z(net_10624) );
CLKBUF_X2 inst_15642 ( .A(net_15489), .Z(net_15490) );
CLKBUF_X2 inst_13091 ( .A(net_12938), .Z(net_12939) );
CLKBUF_X2 inst_10074 ( .A(net_9359), .Z(net_9922) );
NOR2_X1 inst_3620 ( .A2(net_4369), .ZN(net_2001), .A1(net_597) );
CLKBUF_X2 inst_14134 ( .A(net_10998), .Z(net_13982) );
CLKBUF_X2 inst_14763 ( .A(net_10433), .Z(net_14611) );
CLKBUF_X2 inst_9798 ( .A(net_9264), .Z(net_9646) );
XNOR2_X2 inst_260 ( .A(net_2689), .B(net_2671), .ZN(net_1184) );
CLKBUF_X2 inst_11277 ( .A(net_11124), .Z(net_11125) );
CLKBUF_X2 inst_9371 ( .A(net_9218), .Z(net_9219) );
CLKBUF_X2 inst_11597 ( .A(net_11444), .Z(net_11445) );
MUX2_X2 inst_4973 ( .A(net_9023), .Z(net_3937), .B(net_2150), .S(net_622) );
NAND2_X2 inst_4139 ( .ZN(net_5381), .A1(net_5217), .A2(net_5001) );
DFF_X1 inst_6762 ( .Q(net_7542), .D(net_4610), .CK(net_9735) );
NAND2_X2 inst_4611 ( .A2(net_6144), .ZN(net_2619), .A1(net_2618) );
CLKBUF_X2 inst_13839 ( .A(net_13686), .Z(net_13687) );
CLKBUF_X2 inst_10725 ( .A(net_10572), .Z(net_10573) );
NAND2_X2 inst_4567 ( .ZN(net_3083), .A1(net_3082), .A2(net_3081) );
NAND3_X2 inst_3889 ( .ZN(net_5649), .A1(net_5578), .A3(net_5512), .A2(net_5438) );
CLKBUF_X2 inst_17093 ( .A(net_16940), .Z(net_16941) );
CLKBUF_X2 inst_16746 ( .A(net_14432), .Z(net_16594) );
CLKBUF_X2 inst_9880 ( .A(net_9727), .Z(net_9728) );
AOI221_X4 inst_8739 ( .B1(net_8824), .C1(net_8343), .C2(net_6265), .B2(net_6253), .ZN(net_4327), .A(net_4231) );
SDFF_X2 inst_516 ( .Q(net_8870), .D(net_8870), .SI(net_3958), .SE(net_3936), .CK(net_10018) );
CLKBUF_X2 inst_18196 ( .A(net_13416), .Z(net_18044) );
CLKBUF_X2 inst_12243 ( .A(net_12090), .Z(net_12091) );
SDFFR_X2 inst_2258 ( .D(net_7389), .SE(net_2797), .SI(net_198), .Q(net_198), .CK(net_17543), .RN(x6501) );
CLKBUF_X2 inst_13986 ( .A(net_13833), .Z(net_13834) );
XNOR2_X2 inst_190 ( .ZN(net_1594), .B(net_1193), .A(net_1192) );
CLKBUF_X2 inst_16174 ( .A(net_16021), .Z(net_16022) );
CLKBUF_X2 inst_9602 ( .A(net_9377), .Z(net_9450) );
NAND2_X2 inst_4873 ( .A1(net_7480), .A2(net_3921), .ZN(net_1286) );
CLKBUF_X2 inst_13484 ( .A(net_9709), .Z(net_13332) );
CLKBUF_X2 inst_9932 ( .A(net_9471), .Z(net_9780) );
INV_X2 inst_6424 ( .A(net_966), .ZN(net_748) );
SDFFS_X2 inst_2062 ( .SE(net_2417), .SI(net_1330), .Q(net_184), .D(net_184), .CK(net_18103), .SN(x6501) );
CLKBUF_X2 inst_15442 ( .A(net_13446), .Z(net_15290) );
SDFFR_X2 inst_2350 ( .SE(net_2260), .Q(net_315), .D(net_315), .CK(net_11502), .RN(x6501), .SI(x3327) );
CLKBUF_X2 inst_15168 ( .A(net_13493), .Z(net_15016) );
CLKBUF_X2 inst_17471 ( .A(net_17318), .Z(net_17319) );
CLKBUF_X2 inst_15363 ( .A(net_15210), .Z(net_15211) );
CLKBUF_X2 inst_11911 ( .A(net_11758), .Z(net_11759) );
NOR2_X2 inst_3435 ( .A1(net_7651), .A2(net_3081), .ZN(net_3074) );
DFFS_X1 inst_6934 ( .D(net_6145), .CK(net_16347), .SN(x6501), .Q(x890) );
SDFF_X2 inst_829 ( .SI(net_8489), .Q(net_8489), .D(net_3981), .SE(net_3884), .CK(net_12945) );
CLKBUF_X2 inst_15697 ( .A(net_10040), .Z(net_15545) );
XNOR2_X2 inst_197 ( .ZN(net_1547), .B(net_1227), .A(net_1123) );
DFFR_X2 inst_7277 ( .QN(net_7621), .D(net_1842), .CK(net_15668), .RN(x6501) );
NAND2_X2 inst_4702 ( .A1(net_2073), .ZN(net_2050), .A2(net_1784) );
CLKBUF_X2 inst_17628 ( .A(net_17475), .Z(net_17476) );
CLKBUF_X2 inst_10129 ( .A(net_9976), .Z(net_9977) );
CLKBUF_X2 inst_14866 ( .A(net_14713), .Z(net_14714) );
CLKBUF_X2 inst_12830 ( .A(net_12677), .Z(net_12678) );
CLKBUF_X2 inst_17933 ( .A(net_13542), .Z(net_17781) );
CLKBUF_X2 inst_11155 ( .A(net_11002), .Z(net_11003) );
AOI22_X2 inst_8558 ( .A2(net_8250), .B2(net_6117), .A1(net_4800), .ZN(net_2759), .B1(net_2570) );
XNOR2_X2 inst_150 ( .ZN(net_2107), .A(net_1825), .B(net_1824) );
DFF_X1 inst_6743 ( .QN(net_6787), .D(net_5626), .CK(net_11588) );
INV_X4 inst_5358 ( .ZN(net_1147), .A(net_1146) );
NAND2_X2 inst_4540 ( .A2(net_3371), .A1(net_3367), .ZN(net_3366) );
SDFF_X2 inst_887 ( .Q(net_8564), .D(net_8564), .SI(net_3937), .SE(net_3878), .CK(net_12402) );
CLKBUF_X2 inst_18561 ( .A(net_18408), .Z(net_18409) );
CLKBUF_X2 inst_16016 ( .A(net_13055), .Z(net_15864) );
INV_X4 inst_5175 ( .ZN(net_3028), .A(net_2941) );
AOI22_X2 inst_8036 ( .B1(net_8170), .A1(net_7728), .B2(net_6101), .A2(net_6095), .ZN(net_6020) );
CLKBUF_X2 inst_17495 ( .A(net_12243), .Z(net_17343) );
CLKBUF_X2 inst_15630 ( .A(net_11181), .Z(net_15478) );
AOI22_X2 inst_8547 ( .B1(net_6595), .A1(net_6562), .A2(net_6257), .B2(net_6110), .ZN(net_3393) );
CLKBUF_X2 inst_13647 ( .A(net_13494), .Z(net_13495) );
NAND2_X2 inst_4316 ( .A1(net_7057), .A2(net_5162), .ZN(net_5141) );
SDFFR_X2 inst_2357 ( .SE(net_2748), .D(net_2726), .SI(net_473), .Q(net_473), .CK(net_16921), .RN(x6501) );
CLKBUF_X2 inst_13911 ( .A(net_13758), .Z(net_13759) );
INV_X2 inst_6541 ( .A(net_7580), .ZN(net_3139) );
CLKBUF_X2 inst_18180 ( .A(net_18027), .Z(net_18028) );
CLKBUF_X2 inst_12248 ( .A(net_12095), .Z(net_12096) );
SDFF_X2 inst_1961 ( .D(net_7289), .SI(net_6986), .Q(net_6986), .SE(net_6283), .CK(net_15306) );
CLKBUF_X2 inst_14343 ( .A(net_14190), .Z(net_14191) );
INV_X4 inst_5799 ( .A(net_8280), .ZN(net_663) );
INV_X4 inst_5954 ( .A(net_8906), .ZN(net_2786) );
SDFF_X2 inst_1010 ( .SI(net_7322), .Q(net_6663), .D(net_6663), .SE(net_3126), .CK(net_9161) );
AOI22_X2 inst_7934 ( .B1(net_8122), .A1(net_7884), .A2(net_6098), .ZN(net_4191), .B2(net_4190) );
CLKBUF_X2 inst_14939 ( .A(net_10419), .Z(net_14787) );
CLKBUF_X2 inst_14979 ( .A(net_14826), .Z(net_14827) );
SDFF_X2 inst_867 ( .Q(net_8576), .D(net_8576), .SI(net_3957), .SE(net_3878), .CK(net_10971) );
CLKBUF_X2 inst_14179 ( .A(net_14026), .Z(net_14027) );
CLKBUF_X2 inst_18132 ( .A(net_17979), .Z(net_17980) );
NOR2_X2 inst_3568 ( .A2(net_8214), .ZN(net_1456), .A1(net_1175) );
INV_X2 inst_6202 ( .ZN(net_5508), .A(net_5421) );
CLKBUF_X2 inst_16400 ( .A(net_16247), .Z(net_16248) );
CLKBUF_X2 inst_18544 ( .A(net_18391), .Z(net_18392) );
CLKBUF_X2 inst_10760 ( .A(net_10607), .Z(net_10608) );
AOI21_X2 inst_8963 ( .B1(net_6324), .ZN(net_3184), .A(net_3182), .B2(net_3181) );
CLKBUF_X2 inst_15449 ( .A(net_12999), .Z(net_15297) );
CLKBUF_X2 inst_12364 ( .A(net_12211), .Z(net_12212) );
CLKBUF_X2 inst_9342 ( .A(net_9189), .Z(net_9190) );
NAND2_X2 inst_4158 ( .ZN(net_5356), .A2(net_5204), .A1(net_5096) );
CLKBUF_X2 inst_11481 ( .A(net_11328), .Z(net_11329) );
SDFF_X2 inst_1643 ( .SI(net_7717), .Q(net_7717), .D(net_2720), .SE(net_2559), .CK(net_18366) );
NAND2_X2 inst_4660 ( .ZN(net_2415), .A2(net_2315), .A1(net_2314) );
CLKBUF_X2 inst_14537 ( .A(net_11282), .Z(net_14385) );
SDFFR_X2 inst_2120 ( .SI(net_7187), .Q(net_7187), .D(net_6438), .SE(net_4362), .CK(net_17850), .RN(x6501) );
SDFFR_X1 inst_2678 ( .SI(net_7541), .SE(net_5043), .CK(net_9707), .RN(x6501), .Q(x4049), .D(x4049) );
AND2_X2 inst_9196 ( .ZN(net_3386), .A2(net_1727), .A1(net_1507) );
CLKBUF_X2 inst_16898 ( .A(net_16745), .Z(net_16746) );
CLKBUF_X2 inst_15079 ( .A(net_14926), .Z(net_14927) );
SDFFR_X2 inst_2613 ( .Q(net_7381), .D(net_2785), .SE(net_1136), .CK(net_15020), .RN(x6501), .SI(x4707) );
CLKBUF_X2 inst_15003 ( .A(net_11794), .Z(net_14851) );
CLKBUF_X2 inst_10577 ( .A(net_10334), .Z(net_10425) );
DFFR_X2 inst_7143 ( .Q(net_6404), .D(net_2918), .CK(net_18005), .RN(x6501) );
CLKBUF_X2 inst_12239 ( .A(net_9085), .Z(net_12087) );
NAND3_X4 inst_3866 ( .A3(net_6274), .A1(net_6191), .ZN(net_4818), .A2(net_4816) );
CLKBUF_X2 inst_10460 ( .A(net_10307), .Z(net_10308) );
AOI22_X2 inst_8186 ( .B1(net_8679), .A1(net_8642), .B2(net_6109), .A2(net_3857), .ZN(net_3846) );
AOI22_X2 inst_7976 ( .B1(net_8128), .A1(net_7890), .A2(net_6098), .B2(net_4190), .ZN(net_4154) );
CLKBUF_X2 inst_17082 ( .A(net_11410), .Z(net_16930) );
NAND2_X2 inst_4371 ( .A1(net_7154), .A2(net_5166), .ZN(net_5086) );
INV_X4 inst_5253 ( .ZN(net_2282), .A(net_2146) );
CLKBUF_X2 inst_17180 ( .A(net_17027), .Z(net_17028) );
SDFF_X2 inst_1649 ( .SI(net_7730), .Q(net_7730), .D(net_2710), .SE(net_2559), .CK(net_17129) );
AOI22_X2 inst_7756 ( .B1(net_6984), .A1(net_6944), .A2(net_5443), .B2(net_5442), .ZN(net_5382) );
CLKBUF_X2 inst_12921 ( .A(net_10231), .Z(net_12769) );
CLKBUF_X2 inst_13594 ( .A(net_13441), .Z(net_13442) );
INV_X4 inst_5815 ( .A(net_7227), .ZN(net_1612) );
INV_X4 inst_5873 ( .A(net_8283), .ZN(net_975) );
CLKBUF_X2 inst_18557 ( .A(net_15094), .Z(net_18405) );
AOI222_X1 inst_8697 ( .C1(net_7511), .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3200), .B1(net_3136), .A2(net_3008) );
SDFF_X2 inst_669 ( .Q(net_8411), .D(net_8411), .SI(net_3977), .SE(net_3934), .CK(net_10759) );
CLKBUF_X2 inst_9214 ( .A(net_9061), .Z(net_9062) );
CLKBUF_X2 inst_10024 ( .A(net_9224), .Z(net_9872) );
CLKBUF_X2 inst_16092 ( .A(net_15939), .Z(net_15940) );
AOI21_X2 inst_8988 ( .ZN(net_1753), .A(net_1752), .B1(net_1575), .B2(net_1574) );
CLKBUF_X2 inst_14633 ( .A(net_10315), .Z(net_14481) );
CLKBUF_X2 inst_14530 ( .A(net_11530), .Z(net_14378) );
CLKBUF_X2 inst_17817 ( .A(net_17664), .Z(net_17665) );
CLKBUF_X2 inst_10532 ( .A(net_10379), .Z(net_10380) );
AOI22_X2 inst_8236 ( .B1(net_8871), .A1(net_8316), .B2(net_6252), .A2(net_4345), .ZN(net_3801) );
CLKBUF_X2 inst_18056 ( .A(net_13471), .Z(net_17904) );
CLKBUF_X2 inst_17798 ( .A(net_14251), .Z(net_17646) );
NAND2_X2 inst_4897 ( .A2(net_7384), .ZN(net_647), .A1(net_173) );
SDFF_X2 inst_1844 ( .D(net_7288), .SI(net_6945), .Q(net_6945), .SE(net_6281), .CK(net_17682) );
SDFF_X2 inst_1913 ( .D(net_7297), .SI(net_6954), .Q(net_6954), .SE(net_6281), .CK(net_18179) );
INV_X4 inst_5209 ( .A(net_2496), .ZN(net_2382) );
SDFF_X2 inst_1990 ( .SI(net_8052), .Q(net_8052), .D(net_2702), .SE(net_2508), .CK(net_18837) );
INV_X4 inst_5700 ( .A(net_7419), .ZN(net_747) );
XOR2_X2 inst_36 ( .Z(net_1123), .A(net_1122), .B(net_1121) );
CLKBUF_X2 inst_12770 ( .A(net_12617), .Z(net_12618) );
CLKBUF_X2 inst_14658 ( .A(net_14505), .Z(net_14506) );
CLKBUF_X2 inst_13686 ( .A(net_13533), .Z(net_13534) );
AND3_X4 inst_9039 ( .A2(net_6198), .ZN(net_4680), .A1(net_4491), .A3(net_4490) );
CLKBUF_X2 inst_9652 ( .A(net_9409), .Z(net_9500) );
CLKBUF_X2 inst_15175 ( .A(net_12697), .Z(net_15023) );
CLKBUF_X2 inst_18564 ( .A(net_13647), .Z(net_18412) );
CLKBUF_X2 inst_13040 ( .A(net_12887), .Z(net_12888) );
CLKBUF_X2 inst_18011 ( .A(net_13350), .Z(net_17859) );
CLKBUF_X2 inst_16663 ( .A(net_16510), .Z(net_16511) );
CLKBUF_X2 inst_10721 ( .A(net_10568), .Z(net_10569) );
AOI22_X2 inst_7998 ( .B1(net_7927), .A1(net_7825), .B2(net_6103), .A2(net_4398), .ZN(net_4135) );
CLKBUF_X2 inst_19075 ( .A(net_18922), .Z(net_18923) );
AOI22_X2 inst_7954 ( .B1(net_8125), .A1(net_7887), .A2(net_6098), .B2(net_4190), .ZN(net_4173) );
CLKBUF_X2 inst_13284 ( .A(net_13131), .Z(net_13132) );
OAI21_X2 inst_3067 ( .B2(net_6184), .ZN(net_4372), .A(net_4353), .B1(net_1164) );
CLKBUF_X2 inst_13023 ( .A(net_12870), .Z(net_12871) );
CLKBUF_X2 inst_14456 ( .A(net_10566), .Z(net_14304) );
CLKBUF_X2 inst_9877 ( .A(net_9724), .Z(net_9725) );
CLKBUF_X2 inst_17579 ( .A(net_17426), .Z(net_17427) );
AND2_X4 inst_9142 ( .A2(net_5979), .A1(net_5978), .ZN(net_1529) );
CLKBUF_X2 inst_13737 ( .A(net_13584), .Z(net_13585) );
CLKBUF_X2 inst_17572 ( .A(net_17419), .Z(net_17420) );
CLKBUF_X2 inst_10058 ( .A(net_9905), .Z(net_9906) );
INV_X4 inst_5307 ( .ZN(net_1725), .A(net_1098) );
CLKBUF_X2 inst_13188 ( .A(net_9599), .Z(net_13036) );
SDFF_X2 inst_676 ( .Q(net_8703), .D(net_8703), .SI(net_3948), .SE(net_3935), .CK(net_13471) );
CLKBUF_X2 inst_17183 ( .A(net_15655), .Z(net_17031) );
CLKBUF_X2 inst_9755 ( .A(net_9602), .Z(net_9603) );
CLKBUF_X2 inst_16642 ( .A(net_13643), .Z(net_16490) );
CLKBUF_X2 inst_15930 ( .A(net_14388), .Z(net_15778) );
CLKBUF_X2 inst_18660 ( .A(net_18507), .Z(net_18508) );
NAND2_X2 inst_4222 ( .A1(net_7015), .A2(net_5249), .ZN(net_5238) );
HA_X1 inst_6669 ( .S(net_3226), .CO(net_3225), .B(net_3224), .A(net_3192) );
NAND2_X2 inst_4859 ( .ZN(net_2200), .A2(net_864), .A1(net_835) );
CLKBUF_X2 inst_12588 ( .A(net_12435), .Z(net_12436) );
CLKBUF_X2 inst_10193 ( .A(net_9511), .Z(net_10041) );
SDFFR_X2 inst_2255 ( .D(net_7384), .SE(net_2797), .SI(net_193), .Q(net_193), .CK(net_18158), .RN(x6501) );
NAND2_X2 inst_4560 ( .A1(net_3354), .ZN(net_3351), .A2(net_3246) );
SDFF_X2 inst_1076 ( .D(net_7325), .SI(net_6501), .Q(net_6501), .SE(net_3071), .CK(net_11350) );
INV_X2 inst_6360 ( .ZN(net_2168), .A(net_2167) );
INV_X4 inst_6078 ( .A(net_5973), .ZN(x3418) );
CLKBUF_X2 inst_17660 ( .A(net_14400), .Z(net_17508) );
CLKBUF_X2 inst_13292 ( .A(net_12297), .Z(net_13140) );
CLKBUF_X2 inst_9264 ( .A(net_9062), .Z(net_9112) );
SDFF_X2 inst_2000 ( .SI(net_7792), .Q(net_7792), .D(net_2718), .SE(net_2459), .CK(net_18744) );
NAND4_X2 inst_3748 ( .ZN(net_4282), .A1(net_4027), .A2(net_4026), .A3(net_4025), .A4(net_4024) );
DFF_X1 inst_6732 ( .Q(net_6777), .D(net_5637), .CK(net_9208) );
CLKBUF_X2 inst_10223 ( .A(net_9268), .Z(net_10071) );
SDFF_X2 inst_1195 ( .D(net_7317), .SI(net_6526), .Q(net_6526), .SE(net_3086), .CK(net_9824) );
INV_X2 inst_6222 ( .ZN(net_5488), .A(net_5341) );
CLKBUF_X2 inst_16057 ( .A(net_15904), .Z(net_15905) );
CLKBUF_X2 inst_9699 ( .A(net_9546), .Z(net_9547) );
CLKBUF_X2 inst_12252 ( .A(net_12099), .Z(net_12100) );
CLKBUF_X2 inst_11829 ( .A(net_11676), .Z(net_11677) );
DFF_X1 inst_6839 ( .Q(net_6429), .D(net_3608), .CK(net_17978) );
SDFFR_X2 inst_2248 ( .SI(net_7384), .SE(net_2814), .Q(net_243), .D(net_243), .CK(net_17552), .RN(x6501) );
CLKBUF_X2 inst_16740 ( .A(net_16587), .Z(net_16588) );
SDFFR_X2 inst_2453 ( .D(net_7513), .SE(net_2313), .SI(net_429), .Q(net_429), .CK(net_14703), .RN(x6501) );
SDFF_X2 inst_1312 ( .SI(net_7677), .Q(net_7677), .SE(net_2714), .D(net_2658), .CK(net_15544) );
CLKBUF_X2 inst_17166 ( .A(net_17013), .Z(net_17014) );
CLKBUF_X2 inst_18737 ( .A(net_18584), .Z(net_18585) );
CLKBUF_X2 inst_16193 ( .A(net_16040), .Z(net_16041) );
CLKBUF_X2 inst_15145 ( .A(net_11029), .Z(net_14993) );
CLKBUF_X2 inst_18447 ( .A(net_13687), .Z(net_18295) );
INV_X4 inst_5785 ( .A(net_6798), .ZN(net_4355) );
CLKBUF_X2 inst_18141 ( .A(net_17988), .Z(net_17989) );
NOR2_X2 inst_3419 ( .A2(net_7647), .ZN(net_3160), .A1(net_3158) );
CLKBUF_X2 inst_17423 ( .A(net_9812), .Z(net_17271) );
CLKBUF_X2 inst_13749 ( .A(net_13596), .Z(net_13597) );
AOI22_X2 inst_8406 ( .B1(net_8786), .A1(net_8527), .A2(net_3861), .B2(net_3860), .ZN(net_3646) );
MUX2_X2 inst_4951 ( .A(net_7390), .S(net_2378), .Z(net_2373), .B(net_788) );
CLKBUF_X2 inst_14954 ( .A(net_11086), .Z(net_14802) );
CLKBUF_X2 inst_17637 ( .A(net_16342), .Z(net_17485) );
SDFF_X2 inst_971 ( .SI(net_7333), .Q(net_6740), .D(net_6740), .SE(net_3124), .CK(net_9436) );
SDFF_X2 inst_1219 ( .Q(net_7962), .D(net_7962), .SE(net_2755), .SI(net_2718), .CK(net_18825) );
CLKBUF_X2 inst_18246 ( .A(net_12457), .Z(net_18094) );
AOI22_X2 inst_8018 ( .B1(net_8133), .A1(net_7895), .A2(net_6098), .B2(net_4190), .ZN(net_4118) );
NOR2_X2 inst_3459 ( .ZN(net_2874), .A2(net_2747), .A1(net_1469) );
CLKBUF_X2 inst_18345 ( .A(net_18192), .Z(net_18193) );
CLKBUF_X2 inst_16362 ( .A(net_16209), .Z(net_16210) );
NAND2_X2 inst_4488 ( .A2(net_5609), .ZN(net_4484), .A1(net_367) );
CLKBUF_X2 inst_18587 ( .A(net_18434), .Z(net_18435) );
CLKBUF_X2 inst_15357 ( .A(net_15204), .Z(net_15205) );
CLKBUF_X2 inst_12716 ( .A(net_10303), .Z(net_12564) );
CLKBUF_X2 inst_11732 ( .A(net_11579), .Z(net_11580) );
CLKBUF_X2 inst_11741 ( .A(net_10341), .Z(net_11589) );
CLKBUF_X2 inst_15992 ( .A(net_15839), .Z(net_15840) );
CLKBUF_X2 inst_15123 ( .A(net_14970), .Z(net_14971) );
CLKBUF_X2 inst_9454 ( .A(net_9301), .Z(net_9302) );
DFFR_X2 inst_7222 ( .QN(net_7669), .D(net_2259), .CK(net_14579), .RN(x6501) );
CLKBUF_X2 inst_18380 ( .A(net_18227), .Z(net_18228) );
CLKBUF_X2 inst_12628 ( .A(net_10773), .Z(net_12476) );
CLKBUF_X2 inst_12991 ( .A(net_12838), .Z(net_12839) );
CLKBUF_X2 inst_18038 ( .A(net_17885), .Z(net_17886) );
INV_X4 inst_5842 ( .A(net_7382), .ZN(net_978) );
CLKBUF_X2 inst_16206 ( .A(net_16053), .Z(net_16054) );
CLKBUF_X2 inst_10135 ( .A(net_9982), .Z(net_9983) );
NOR3_X2 inst_3286 ( .ZN(net_2311), .A3(net_2310), .A2(net_2234), .A1(net_1737) );
NAND2_X2 inst_4225 ( .A1(net_6896), .A2(net_5247), .ZN(net_5235) );
INV_X4 inst_5625 ( .A(net_6462), .ZN(net_1667) );
CLKBUF_X2 inst_11371 ( .A(net_11218), .Z(net_11219) );
CLKBUF_X2 inst_11421 ( .A(net_11268), .Z(net_11269) );
CLKBUF_X2 inst_9533 ( .A(net_9287), .Z(net_9381) );
NAND2_X2 inst_4141 ( .ZN(net_5379), .A2(net_5216), .A1(net_5114) );
CLKBUF_X2 inst_14293 ( .A(net_14140), .Z(net_14141) );
NAND2_X2 inst_4591 ( .A1(net_8254), .A2(net_6100), .ZN(net_3022) );
CLKBUF_X2 inst_16470 ( .A(net_16317), .Z(net_16318) );
INV_X4 inst_5318 ( .ZN(net_1586), .A(net_1454) );
CLKBUF_X2 inst_12493 ( .A(net_12340), .Z(net_12341) );
CLKBUF_X2 inst_9865 ( .A(net_9226), .Z(net_9713) );
CLKBUF_X2 inst_17119 ( .A(net_16966), .Z(net_16967) );
AND2_X2 inst_9162 ( .ZN(net_2831), .A1(net_2754), .A2(net_2753) );
CLKBUF_X2 inst_11290 ( .A(net_11137), .Z(net_11138) );
XNOR2_X2 inst_188 ( .A(net_1792), .B(net_1788), .ZN(net_1640) );
NAND2_X2 inst_4528 ( .A2(net_3566), .ZN(net_3558), .A1(net_3557) );
CLKBUF_X2 inst_13534 ( .A(net_13381), .Z(net_13382) );
INV_X4 inst_6093 ( .A(net_8948), .ZN(net_658) );
CLKBUF_X2 inst_14586 ( .A(net_14433), .Z(net_14434) );
CLKBUF_X2 inst_18732 ( .A(net_18579), .Z(net_18580) );
OAI21_X2 inst_3011 ( .ZN(net_5719), .A(net_5718), .B2(net_5587), .B1(net_4823) );
CLKBUF_X2 inst_18761 ( .A(net_12856), .Z(net_18609) );
CLKBUF_X2 inst_16585 ( .A(net_16432), .Z(net_16433) );
NAND2_X2 inst_4826 ( .A2(net_5957), .ZN(net_1107), .A1(net_1106) );
HA_X1 inst_6695 ( .S(net_2822), .CO(net_2821), .B(net_2505), .A(x3079) );
SDFF_X2 inst_1537 ( .Q(net_7990), .D(net_7990), .SI(net_2589), .SE(net_2542), .CK(net_18865) );
SDFF_X2 inst_2041 ( .SI(net_7790), .Q(net_7790), .D(net_2590), .SE(net_2459), .CK(net_15943) );
INV_X2 inst_6323 ( .ZN(net_3340), .A(net_3283) );
INV_X4 inst_5235 ( .ZN(net_2260), .A(net_2196) );
CLKBUF_X2 inst_15509 ( .A(net_15189), .Z(net_15357) );
NAND2_X2 inst_4589 ( .ZN(net_2882), .A2(net_2881), .A1(net_1446) );
DFF_X1 inst_6768 ( .Q(net_7547), .D(net_4604), .CK(net_9719) );
CLKBUF_X2 inst_18443 ( .A(net_11357), .Z(net_18291) );
CLKBUF_X2 inst_11550 ( .A(net_9219), .Z(net_11398) );
NOR2_X4 inst_3325 ( .ZN(net_3598), .A2(net_3597), .A1(net_3251) );
CLKBUF_X2 inst_13393 ( .A(net_13240), .Z(net_13241) );
CLKBUF_X2 inst_11145 ( .A(net_10992), .Z(net_10993) );
CLKBUF_X2 inst_11085 ( .A(net_10932), .Z(net_10933) );
AND2_X4 inst_9083 ( .ZN(net_2889), .A2(net_2888), .A1(net_2528) );
CLKBUF_X2 inst_13991 ( .A(net_11762), .Z(net_13839) );
NAND2_X2 inst_4168 ( .ZN(net_5343), .A2(net_5198), .A1(net_5087) );
XNOR2_X2 inst_195 ( .A(net_7660), .ZN(net_1550), .B(net_1549) );
CLKBUF_X2 inst_18507 ( .A(net_18354), .Z(net_18355) );
CLKBUF_X2 inst_11835 ( .A(net_10378), .Z(net_11683) );
CLKBUF_X2 inst_12839 ( .A(net_12686), .Z(net_12687) );
SDFF_X2 inst_1987 ( .D(net_7288), .SI(net_6905), .Q(net_6905), .SE(net_6284), .CK(net_14869) );
CLKBUF_X2 inst_13418 ( .A(net_13265), .Z(net_13266) );
CLKBUF_X2 inst_14372 ( .A(net_9154), .Z(net_14220) );
INV_X4 inst_5605 ( .A(net_9055), .ZN(net_2827) );
DFFR_X2 inst_7070 ( .QN(net_7418), .D(net_4201), .CK(net_12301), .RN(x6501) );
DFFR_X2 inst_7106 ( .QN(net_6329), .D(net_3209), .CK(net_14728), .RN(x6501) );
NAND2_X2 inst_4780 ( .ZN(net_1701), .A2(net_1129), .A1(net_1104) );
CLKBUF_X2 inst_12981 ( .A(net_12828), .Z(net_12829) );
CLKBUF_X2 inst_15468 ( .A(net_15315), .Z(net_15316) );
NAND2_X2 inst_4658 ( .A1(net_2735), .A2(net_2334), .ZN(net_2270) );
INV_X4 inst_5916 ( .ZN(net_2733), .A(net_271) );
DFFR_X2 inst_7154 ( .QN(net_9051), .D(net_2851), .CK(net_11157), .RN(x6501) );
SDFF_X2 inst_1589 ( .Q(net_8016), .D(net_8016), .SI(net_2708), .SE(net_2545), .CK(net_15521) );
CLKBUF_X2 inst_11994 ( .A(net_9739), .Z(net_11842) );
AOI21_X2 inst_8926 ( .B2(net_5871), .ZN(net_5687), .A(net_5677), .B1(net_2750) );
CLKBUF_X2 inst_14114 ( .A(net_13961), .Z(net_13962) );
INV_X4 inst_5607 ( .A(net_6824), .ZN(net_1029) );
CLKBUF_X2 inst_14095 ( .A(net_13942), .Z(net_13943) );
CLKBUF_X2 inst_16499 ( .A(net_16346), .Z(net_16347) );
CLKBUF_X2 inst_15263 ( .A(net_9587), .Z(net_15111) );
CLKBUF_X2 inst_15160 ( .A(net_15007), .Z(net_15008) );
XNOR2_X2 inst_335 ( .B(net_7379), .A(net_6361), .ZN(net_792) );
CLKBUF_X2 inst_15244 ( .A(net_15091), .Z(net_15092) );
CLKBUF_X2 inst_12827 ( .A(net_12674), .Z(net_12675) );
CLKBUF_X2 inst_14406 ( .A(net_14253), .Z(net_14254) );
DFFS_X2 inst_6862 ( .QN(net_6332), .D(net_5581), .CK(net_18939), .SN(x6501) );
AOI22_X2 inst_8420 ( .B1(net_6520), .A1(net_6487), .A2(net_6137), .B2(net_6104), .ZN(net_3522) );
CLKBUF_X2 inst_9336 ( .A(net_9183), .Z(net_9184) );
CLKBUF_X2 inst_11562 ( .A(net_9273), .Z(net_11410) );
CLKBUF_X2 inst_14045 ( .A(net_13892), .Z(net_13893) );
CLKBUF_X2 inst_16155 ( .A(net_9060), .Z(net_16003) );
CLKBUF_X2 inst_14276 ( .A(net_9264), .Z(net_14124) );
SDFF_X2 inst_438 ( .Q(net_8766), .D(net_8766), .SE(net_3982), .SI(net_3954), .CK(net_12639) );
CLKBUF_X2 inst_13311 ( .A(net_10201), .Z(net_13159) );
DFFR_X2 inst_7326 ( .QN(net_400), .D(net_398), .CK(net_11605), .RN(x6501) );
INV_X2 inst_6351 ( .ZN(net_2286), .A(net_2215) );
CLKBUF_X2 inst_10769 ( .A(net_10616), .Z(net_10617) );
CLKBUF_X2 inst_14336 ( .A(net_13043), .Z(net_14184) );
CLKBUF_X2 inst_9692 ( .A(net_9539), .Z(net_9540) );
XNOR2_X2 inst_324 ( .B(net_7368), .ZN(net_935), .A(net_493) );
CLKBUF_X2 inst_11640 ( .A(net_11487), .Z(net_11488) );
NOR2_X2 inst_3550 ( .A1(net_1925), .ZN(net_1900), .A2(net_1475) );
INV_X4 inst_6046 ( .A(net_6308), .ZN(net_2682) );
NAND2_X2 inst_4083 ( .ZN(net_5852), .A2(net_5751), .A1(net_549) );
CLKBUF_X2 inst_17240 ( .A(net_17087), .Z(net_17088) );
XOR2_X2 inst_43 ( .A(net_6204), .Z(net_1042), .B(net_554) );
INV_X4 inst_5936 ( .A(net_7246), .ZN(net_1867) );
SDFF_X2 inst_1707 ( .SI(net_7852), .Q(net_7852), .D(net_2574), .SE(net_2558), .CK(net_16027) );
CLKBUF_X2 inst_17955 ( .A(net_17337), .Z(net_17803) );
DFFR_X2 inst_7213 ( .D(net_2379), .QN(net_229), .CK(net_14786), .RN(x6501) );
DFF_X1 inst_6715 ( .QN(net_6791), .D(net_5622), .CK(net_11601) );
AOI22_X2 inst_8115 ( .B1(net_8047), .A1(net_7843), .B2(net_6107), .A2(net_4400), .ZN(net_4033) );
SDFF_X2 inst_375 ( .SI(net_8309), .Q(net_8309), .SE(net_3978), .D(net_3945), .CK(net_13372) );
CLKBUF_X2 inst_11241 ( .A(net_10501), .Z(net_11089) );
CLKBUF_X2 inst_9959 ( .A(net_9806), .Z(net_9807) );
AOI222_X1 inst_8606 ( .B2(net_6778), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5818), .A1(net_3218), .C1(x2633) );
NOR2_X2 inst_3490 ( .A1(net_7299), .ZN(net_2433), .A2(net_2146) );
DFFR_X2 inst_7039 ( .QN(net_7510), .D(net_4845), .CK(net_14840), .RN(x6501) );
CLKBUF_X2 inst_15780 ( .A(net_11906), .Z(net_15628) );
CLKBUF_X2 inst_10933 ( .A(net_10780), .Z(net_10781) );
XNOR2_X2 inst_285 ( .A(net_6836), .B(net_1029), .ZN(net_1010) );
DFFR_X2 inst_7215 ( .D(net_2375), .QN(net_230), .CK(net_15001), .RN(x6501) );
SDFF_X2 inst_1830 ( .D(net_7292), .SI(net_6869), .Q(net_6869), .SE(net_6282), .CK(net_14895) );
CLKBUF_X2 inst_18515 ( .A(net_18362), .Z(net_18363) );
CLKBUF_X2 inst_11780 ( .A(net_10674), .Z(net_11628) );
INV_X4 inst_5563 ( .A(net_845), .ZN(net_604) );
SDFF_X2 inst_1563 ( .Q(net_8010), .D(net_8010), .SI(net_2721), .SE(net_2545), .CK(net_15770) );
INV_X2 inst_6363 ( .A(net_4385), .ZN(net_2106) );
CLKBUF_X2 inst_17044 ( .A(net_16891), .Z(net_16892) );
NOR4_X2 inst_3242 ( .ZN(net_1626), .A1(net_1625), .A2(net_1236), .A3(net_868), .A4(net_857) );
DFFR_X1 inst_7398 ( .D(net_5760), .CK(net_16773), .RN(x6501), .Q(x480) );
CLKBUF_X2 inst_10638 ( .A(net_10485), .Z(net_10486) );
CLKBUF_X2 inst_9895 ( .A(net_9657), .Z(net_9743) );
SDFF_X2 inst_982 ( .SI(net_7318), .Q(net_6725), .D(net_6725), .SE(net_3124), .CK(net_12122) );
OAI21_X2 inst_3138 ( .ZN(net_2061), .B2(net_2060), .A(net_2050), .B1(net_729) );
CLKBUF_X2 inst_17451 ( .A(net_16436), .Z(net_17299) );
CLKBUF_X2 inst_10864 ( .A(net_10711), .Z(net_10712) );
XNOR2_X2 inst_299 ( .B(net_1118), .ZN(net_983), .A(net_598) );
CLKBUF_X2 inst_13871 ( .A(net_13718), .Z(net_13719) );
CLKBUF_X2 inst_10567 ( .A(net_10414), .Z(net_10415) );
SDFF_X2 inst_1798 ( .D(net_7280), .SI(net_6977), .Q(net_6977), .SE(net_6283), .CK(net_19011) );
OAI22_X2 inst_2927 ( .B1(net_9054), .A2(net_2963), .ZN(net_2854), .B2(net_2852), .A1(net_1920) );
CLKBUF_X2 inst_10336 ( .A(net_10183), .Z(net_10184) );
INV_X4 inst_5853 ( .A(net_6348), .ZN(net_2137) );
CLKBUF_X2 inst_10383 ( .A(net_10230), .Z(net_10231) );
CLKBUF_X2 inst_17826 ( .A(net_14723), .Z(net_17674) );
CLKBUF_X2 inst_17016 ( .A(net_16863), .Z(net_16864) );
AOI221_X4 inst_8727 ( .B1(net_8842), .C1(net_8361), .C2(net_6265), .B2(net_6253), .ZN(net_4338), .A(net_4248) );
SDFFR_X1 inst_2760 ( .SI(net_7595), .Q(net_7595), .SE(net_3144), .D(net_1506), .CK(net_13457), .RN(x6501) );
INV_X2 inst_6452 ( .A(net_6420), .ZN(net_590) );
CLKBUF_X2 inst_18838 ( .A(net_18685), .Z(net_18686) );
CLKBUF_X2 inst_15213 ( .A(net_15060), .Z(net_15061) );
DFFR_X2 inst_7098 ( .QN(net_6470), .D(net_3344), .CK(net_15101), .RN(x6501) );
CLKBUF_X2 inst_17596 ( .A(net_17443), .Z(net_17444) );
INV_X2 inst_6288 ( .ZN(net_4211), .A(net_3919) );
DFFR_X2 inst_7030 ( .QN(net_7488), .D(net_5046), .CK(net_16683), .RN(x6501) );
CLKBUF_X2 inst_15581 ( .A(net_15428), .Z(net_15429) );
INV_X4 inst_5129 ( .ZN(net_4402), .A(net_4354) );
CLKBUF_X2 inst_13524 ( .A(net_13371), .Z(net_13372) );
CLKBUF_X2 inst_14841 ( .A(net_14688), .Z(net_14689) );
CLKBUF_X2 inst_10656 ( .A(net_10503), .Z(net_10504) );
MUX2_X2 inst_4995 ( .A(net_9040), .Z(net_3954), .B(net_3390), .S(net_622) );
NOR3_X2 inst_3260 ( .A3(net_4513), .ZN(net_3322), .A1(net_3191), .A2(net_2643) );
OAI21_X2 inst_3158 ( .B2(net_2048), .ZN(net_1971), .A(net_1970), .B1(net_1690) );
NAND2_X2 inst_4190 ( .ZN(net_5310), .A1(net_5183), .A2(net_4984) );
CLKBUF_X2 inst_17878 ( .A(net_9729), .Z(net_17726) );
CLKBUF_X2 inst_13894 ( .A(net_11859), .Z(net_13742) );
CLKBUF_X2 inst_11248 ( .A(net_9414), .Z(net_11096) );
INV_X4 inst_5387 ( .A(net_7209), .ZN(net_1327) );
CLKBUF_X2 inst_14067 ( .A(net_13914), .Z(net_13915) );
SDFFR_X2 inst_2186 ( .QN(net_9005), .SE(net_2776), .D(net_2774), .SI(net_2529), .CK(net_18909), .RN(x6501) );
NOR3_X2 inst_3269 ( .A1(net_6126), .ZN(net_2533), .A2(net_2532), .A3(net_2531) );
CLKBUF_X2 inst_15745 ( .A(net_15592), .Z(net_15593) );
SDFF_X2 inst_1944 ( .SI(net_8047), .Q(net_8047), .D(net_2655), .SE(net_2508), .CK(net_18515) );
AND2_X4 inst_9079 ( .ZN(net_3124), .A2(net_2940), .A1(net_2904) );
XNOR2_X2 inst_210 ( .B(net_8896), .A(net_3363), .ZN(net_1464) );
CLKBUF_X2 inst_13763 ( .A(net_13610), .Z(net_13611) );
CLKBUF_X2 inst_11675 ( .A(net_11522), .Z(net_11523) );
OAI21_X2 inst_3101 ( .ZN(net_2653), .B1(net_2652), .B2(net_2428), .A(net_1837) );
CLKBUF_X2 inst_16142 ( .A(net_15989), .Z(net_15990) );
MUX2_X2 inst_4942 ( .B(net_6318), .S(net_5522), .Z(net_2638), .A(net_2637) );
CLKBUF_X2 inst_14998 ( .A(net_14845), .Z(net_14846) );
INV_X4 inst_5331 ( .ZN(net_2389), .A(net_1346) );
AOI22_X2 inst_8164 ( .B1(net_8741), .A1(net_8371), .ZN(net_3871), .A2(net_3867), .B2(net_3866) );
DFFR_X2 inst_7123 ( .Q(net_8257), .D(net_3180), .CK(net_18495), .RN(x6501) );
SDFF_X2 inst_1294 ( .Q(net_7816), .D(net_7816), .SE(net_2730), .SI(net_2584), .CK(net_15632) );
CLKBUF_X2 inst_16865 ( .A(net_16712), .Z(net_16713) );
SDFF_X2 inst_1712 ( .Q(net_7903), .D(net_7903), .SI(net_2660), .SE(net_2543), .CK(net_14257) );
INV_X4 inst_5238 ( .ZN(net_2334), .A(net_2013) );
CLKBUF_X2 inst_14605 ( .A(net_14452), .Z(net_14453) );
OAI21_X2 inst_3108 ( .B2(net_2489), .ZN(net_2484), .A(net_2335), .B1(net_1758) );
CLKBUF_X2 inst_12626 ( .A(net_12473), .Z(net_12474) );
OR2_X4 inst_2853 ( .A1(net_7401), .ZN(net_1380), .A2(net_656) );
DFFR_X2 inst_7267 ( .QN(net_6381), .D(net_1993), .CK(net_15928), .RN(x6501) );
CLKBUF_X2 inst_15331 ( .A(net_15178), .Z(net_15179) );
CLKBUF_X2 inst_10291 ( .A(net_10138), .Z(net_10139) );
INV_X2 inst_6546 ( .A(net_6474), .ZN(net_3282) );
CLKBUF_X2 inst_12166 ( .A(net_12013), .Z(net_12014) );
AOI22_X2 inst_7855 ( .A2(net_5595), .ZN(net_4652), .B2(net_4388), .B1(net_2606), .A1(net_326) );
CLKBUF_X2 inst_15055 ( .A(net_14902), .Z(net_14903) );
AOI22_X2 inst_8553 ( .B2(net_4889), .A1(net_4803), .ZN(net_3057), .B1(net_3056), .A2(net_2927) );
CLKBUF_X2 inst_11658 ( .A(net_11505), .Z(net_11506) );
CLKBUF_X2 inst_10853 ( .A(net_10700), .Z(net_10701) );
CLKBUF_X2 inst_18651 ( .A(net_18498), .Z(net_18499) );
INV_X2 inst_6291 ( .ZN(net_4207), .A(net_3916) );
CLKBUF_X2 inst_14848 ( .A(net_11582), .Z(net_14696) );
CLKBUF_X2 inst_12476 ( .A(net_12323), .Z(net_12324) );
CLKBUF_X2 inst_14547 ( .A(net_14394), .Z(net_14395) );
INV_X4 inst_5740 ( .A(net_6414), .ZN(net_564) );
CLKBUF_X2 inst_10602 ( .A(net_10449), .Z(net_10450) );
CLKBUF_X2 inst_10993 ( .A(net_10481), .Z(net_10841) );
INV_X2 inst_6227 ( .ZN(net_5483), .A(net_5318) );
CLKBUF_X2 inst_13489 ( .A(net_13336), .Z(net_13337) );
CLKBUF_X2 inst_14930 ( .A(net_14777), .Z(net_14778) );
CLKBUF_X2 inst_15511 ( .A(net_15358), .Z(net_15359) );
CLKBUF_X2 inst_18613 ( .A(net_18460), .Z(net_18461) );
CLKBUF_X2 inst_14898 ( .A(net_12017), .Z(net_14746) );
CLKBUF_X2 inst_11620 ( .A(net_11467), .Z(net_11468) );
CLKBUF_X2 inst_11605 ( .A(net_11452), .Z(net_11453) );
SDFF_X2 inst_907 ( .SI(net_8725), .Q(net_8725), .SE(net_6195), .D(net_3956), .CK(net_10051) );
SDFF_X2 inst_922 ( .SI(net_8710), .Q(net_8710), .SE(net_6195), .D(net_3947), .CK(net_12400) );
CLKBUF_X2 inst_11323 ( .A(net_11170), .Z(net_11171) );
CLKBUF_X2 inst_18095 ( .A(net_10520), .Z(net_17943) );
AOI22_X2 inst_8225 ( .B1(net_8796), .A1(net_8537), .A2(net_3861), .B2(net_3860), .ZN(net_3812) );
CLKBUF_X2 inst_18387 ( .A(net_12670), .Z(net_18235) );
AOI221_X2 inst_8773 ( .B1(net_5268), .C2(net_5267), .ZN(net_5266), .A(net_4916), .B2(net_4636), .C1(net_177) );
CLKBUF_X2 inst_19111 ( .A(net_18958), .Z(net_18959) );
CLKBUF_X2 inst_15072 ( .A(net_11094), .Z(net_14920) );
CLKBUF_X2 inst_12435 ( .A(net_12282), .Z(net_12283) );
CLKBUF_X2 inst_10693 ( .A(net_10540), .Z(net_10541) );
CLKBUF_X2 inst_9475 ( .A(net_9322), .Z(net_9323) );
CLKBUF_X2 inst_14418 ( .A(net_14265), .Z(net_14266) );
AOI22_X2 inst_8516 ( .B1(net_6551), .A1(net_6518), .A2(net_6137), .B2(net_6104), .ZN(net_3424) );
CLKBUF_X2 inst_12621 ( .A(net_12468), .Z(net_12469) );
CLKBUF_X2 inst_13231 ( .A(net_10877), .Z(net_13079) );
NAND3_X2 inst_3907 ( .ZN(net_5631), .A1(net_5560), .A3(net_5494), .A2(net_5366) );
CLKBUF_X2 inst_9619 ( .A(net_9466), .Z(net_9467) );
CLKBUF_X2 inst_14752 ( .A(net_9329), .Z(net_14600) );
CLKBUF_X2 inst_12383 ( .A(net_12230), .Z(net_12231) );
NAND4_X2 inst_3692 ( .A4(net_6248), .A1(net_6247), .ZN(net_4445), .A2(net_3813), .A3(net_3812) );
CLKBUF_X2 inst_18033 ( .A(net_17880), .Z(net_17881) );
SDFF_X2 inst_653 ( .Q(net_8425), .D(net_8425), .SI(net_3967), .SE(net_3934), .CK(net_13040) );
AOI22_X2 inst_8304 ( .A1(net_8621), .B1(net_8436), .A2(net_3864), .B2(net_3863), .ZN(net_3741) );
SDFF_X2 inst_1746 ( .SI(net_7301), .Q(net_7158), .D(net_7158), .SE(net_6279), .CK(net_15893) );
CLKBUF_X2 inst_11099 ( .A(net_10946), .Z(net_10947) );
CLKBUF_X2 inst_18274 ( .A(net_11063), .Z(net_18122) );
CLKBUF_X2 inst_13406 ( .A(net_13253), .Z(net_13254) );
AOI22_X2 inst_8233 ( .B1(net_8797), .A1(net_8538), .A2(net_3861), .B2(net_3860), .ZN(net_3804) );
CLKBUF_X2 inst_15817 ( .A(net_13282), .Z(net_15665) );
NAND4_X2 inst_3649 ( .A4(net_5996), .A1(net_5995), .ZN(net_4616), .A2(net_4199), .A3(net_4198) );
CLKBUF_X2 inst_17131 ( .A(net_16978), .Z(net_16979) );
NAND2_X2 inst_4609 ( .A2(net_6144), .ZN(net_2623), .A1(net_2622) );
INV_X2 inst_6526 ( .A(net_7669), .ZN(net_526) );
CLKBUF_X2 inst_11843 ( .A(net_11445), .Z(net_11691) );
SDFFR_X1 inst_2656 ( .D(net_6778), .SE(net_4506), .CK(net_11418), .RN(x6501), .SI(x1532), .Q(x1532) );
CLKBUF_X2 inst_16165 ( .A(net_10826), .Z(net_16013) );
AOI22_X2 inst_8301 ( .B1(net_8732), .A1(net_8510), .ZN(net_6069), .B2(net_4350), .A2(net_4349) );
SDFF_X2 inst_1604 ( .Q(net_8140), .D(net_8140), .SI(net_2715), .SE(net_2541), .CK(net_14164) );
CLKBUF_X2 inst_18146 ( .A(net_17993), .Z(net_17994) );
CLKBUF_X2 inst_9426 ( .A(net_9180), .Z(net_9274) );
CLKBUF_X2 inst_18818 ( .A(net_18665), .Z(net_18666) );
CLKBUF_X2 inst_13854 ( .A(net_12068), .Z(net_13702) );
CLKBUF_X2 inst_14441 ( .A(net_10617), .Z(net_14289) );
AOI222_X2 inst_8592 ( .C1(net_7516), .A1(net_6177), .C2(net_4889), .B2(net_4888), .A2(net_4803), .ZN(net_3874), .B1(net_3134) );
CLKBUF_X2 inst_16934 ( .A(net_11120), .Z(net_16782) );
XOR2_X2 inst_7 ( .Z(net_2507), .A(net_2496), .B(net_2493) );
CLKBUF_X2 inst_18642 ( .A(net_18489), .Z(net_18490) );
CLKBUF_X2 inst_9672 ( .A(net_9519), .Z(net_9520) );
CLKBUF_X2 inst_16465 ( .A(net_16312), .Z(net_16313) );
NOR2_X2 inst_3450 ( .ZN(net_2980), .A2(net_2973), .A1(net_1345) );
CLKBUF_X2 inst_9707 ( .A(net_9554), .Z(net_9555) );
CLKBUF_X2 inst_13742 ( .A(net_13589), .Z(net_13590) );
INV_X4 inst_5408 ( .ZN(net_1095), .A(net_875) );
CLKBUF_X2 inst_17074 ( .A(net_11013), .Z(net_16922) );
CLKBUF_X2 inst_12036 ( .A(net_10494), .Z(net_11884) );
SDFF_X2 inst_1136 ( .D(net_7314), .SI(net_6556), .Q(net_6556), .SE(net_3070), .CK(net_9916) );
CLKBUF_X2 inst_10402 ( .A(net_10249), .Z(net_10250) );
CLKBUF_X2 inst_13360 ( .A(net_13207), .Z(net_13208) );
CLKBUF_X2 inst_11262 ( .A(net_11109), .Z(net_11110) );
CLKBUF_X2 inst_19069 ( .A(net_14372), .Z(net_18917) );
CLKBUF_X2 inst_16141 ( .A(net_15988), .Z(net_15989) );
CLKBUF_X2 inst_9621 ( .A(net_9407), .Z(net_9469) );
CLKBUF_X2 inst_14474 ( .A(net_14321), .Z(net_14322) );
NOR3_X2 inst_3311 ( .A2(net_7221), .A1(net_3162), .ZN(net_1733), .A3(net_1520) );
CLKBUF_X2 inst_13598 ( .A(net_13445), .Z(net_13446) );
CLKBUF_X2 inst_13339 ( .A(net_12910), .Z(net_13187) );
INV_X4 inst_5081 ( .ZN(net_5754), .A(net_5722) );
INV_X4 inst_5117 ( .A(net_8224), .ZN(net_4849) );
MUX2_X2 inst_4929 ( .Z(net_3261), .A(net_3219), .B(net_3018), .S(x3685) );
INV_X4 inst_5114 ( .ZN(net_4973), .A(x1130) );
CLKBUF_X2 inst_13942 ( .A(net_10403), .Z(net_13790) );
CLKBUF_X2 inst_14885 ( .A(net_14732), .Z(net_14733) );
CLKBUF_X2 inst_10423 ( .A(net_9335), .Z(net_10271) );
DFFR_X2 inst_7341 ( .Q(net_7331), .CK(net_11664), .D(x13004), .RN(x6501) );
INV_X2 inst_6268 ( .A(net_8227), .ZN(net_4629) );
CLKBUF_X2 inst_17753 ( .A(net_10996), .Z(net_17601) );
NAND4_X2 inst_3713 ( .ZN(net_4424), .A4(net_4331), .A1(net_3680), .A2(net_3679), .A3(net_3678) );
INV_X4 inst_5681 ( .ZN(net_576), .A(net_276) );
SDFFR_X2 inst_2394 ( .SE(net_2260), .Q(net_314), .D(net_314), .CK(net_10455), .RN(x6501), .SI(x3372) );
NAND2_X2 inst_4574 ( .A1(net_8261), .A2(net_2996), .ZN(net_2995) );
AOI22_X2 inst_8562 ( .A1(net_2699), .A2(net_2334), .B2(net_2333), .ZN(net_2332), .B1(net_2039) );
CLKBUF_X2 inst_9404 ( .A(net_9130), .Z(net_9252) );
CLKBUF_X2 inst_10681 ( .A(net_10528), .Z(net_10529) );
CLKBUF_X2 inst_10612 ( .A(net_10459), .Z(net_10460) );
INV_X4 inst_5294 ( .A(net_1814), .ZN(net_1688) );
CLKBUF_X2 inst_17962 ( .A(net_17809), .Z(net_17810) );
INV_X4 inst_5251 ( .A(net_2127), .ZN(net_1857) );
NAND2_X2 inst_4422 ( .A1(net_6860), .A2(net_5016), .ZN(net_5005) );
CLKBUF_X2 inst_12578 ( .A(net_12425), .Z(net_12426) );
CLKBUF_X2 inst_12219 ( .A(net_11819), .Z(net_12067) );
CLKBUF_X2 inst_14056 ( .A(net_13903), .Z(net_13904) );
CLKBUF_X2 inst_11905 ( .A(net_11752), .Z(net_11753) );
AOI222_X1 inst_8623 ( .A2(net_8228), .B2(net_5535), .A1(net_5268), .ZN(net_4882), .C2(net_4881), .B1(net_454), .C1(net_235) );
INV_X4 inst_5092 ( .ZN(net_5705), .A(net_5681) );
CLKBUF_X2 inst_15330 ( .A(net_15177), .Z(net_15178) );
INV_X4 inst_5342 ( .A(net_1836), .ZN(net_1379) );
SDFF_X2 inst_1670 ( .SI(net_7769), .Q(net_7769), .D(net_2716), .SE(net_2560), .CK(net_17063) );
CLKBUF_X2 inst_12932 ( .A(net_9353), .Z(net_12780) );
CLKBUF_X2 inst_11491 ( .A(net_11338), .Z(net_11339) );
CLKBUF_X2 inst_10352 ( .A(net_9986), .Z(net_10200) );
AOI222_X1 inst_8646 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3920), .B1(net_3016), .C1(net_3014), .A1(x13826) );
AND4_X4 inst_9028 ( .ZN(net_2974), .A2(net_2868), .A1(net_1443), .A3(net_556), .A4(net_541) );
CLKBUF_X2 inst_16512 ( .A(net_13970), .Z(net_16360) );
CLKBUF_X2 inst_10677 ( .A(net_10524), .Z(net_10525) );
CLKBUF_X2 inst_10327 ( .A(net_10131), .Z(net_10175) );
INV_X8 inst_5027 ( .ZN(net_3880), .A(net_3306) );
INV_X4 inst_5883 ( .A(net_8893), .ZN(net_1167) );
OAI21_X2 inst_3113 ( .ZN(net_2434), .B2(net_2433), .A(net_2431), .B1(net_1147) );
CLKBUF_X2 inst_13500 ( .A(net_13347), .Z(net_13348) );
CLKBUF_X2 inst_19074 ( .A(net_18921), .Z(net_18922) );
CLKBUF_X2 inst_18775 ( .A(net_18622), .Z(net_18623) );
NAND4_X2 inst_3695 ( .ZN(net_4442), .A4(net_4342), .A1(net_3793), .A2(net_3792), .A3(net_3791) );
CLKBUF_X2 inst_12309 ( .A(net_12156), .Z(net_12157) );
HA_X1 inst_6687 ( .S(net_2979), .CO(net_2978), .B(net_2874), .A(x2805) );
SDFFR_X2 inst_2385 ( .SE(net_2260), .Q(net_372), .D(net_372), .CK(net_11456), .RN(x6501), .SI(x1597) );
SDFFR_X2 inst_2336 ( .D(net_7367), .SE(net_2738), .SI(net_1914), .QN(net_263), .CK(net_13551), .RN(x6501) );
CLKBUF_X2 inst_18061 ( .A(net_13401), .Z(net_17909) );
CLKBUF_X2 inst_16044 ( .A(net_15891), .Z(net_15892) );
INV_X4 inst_5927 ( .ZN(net_2693), .A(net_279) );
AOI22_X2 inst_8574 ( .A1(net_2547), .B2(net_1919), .A2(net_1918), .ZN(net_1915), .B1(net_1914) );
CLKBUF_X2 inst_13549 ( .A(net_13396), .Z(net_13397) );
CLKBUF_X2 inst_9482 ( .A(net_9288), .Z(net_9330) );
CLKBUF_X2 inst_17263 ( .A(net_17110), .Z(net_17111) );
XNOR2_X2 inst_223 ( .ZN(net_1388), .B(net_1387), .A(net_620) );
DFF_X1 inst_6814 ( .Q(net_8228), .D(net_4453), .CK(net_17219) );
INV_X4 inst_5278 ( .ZN(net_1684), .A(net_1461) );
INV_X4 inst_6042 ( .A(net_7358), .ZN(net_665) );
CLKBUF_X2 inst_15884 ( .A(net_15731), .Z(net_15732) );
CLKBUF_X2 inst_13811 ( .A(net_9962), .Z(net_13659) );
SDFFR_X2 inst_2420 ( .D(net_2682), .SE(net_2313), .SI(net_467), .Q(net_467), .CK(net_17450), .RN(x6501) );
NOR2_X2 inst_3564 ( .A1(net_1655), .ZN(net_1287), .A2(net_1286) );
CLKBUF_X2 inst_19150 ( .A(net_18997), .Z(net_18998) );
CLKBUF_X2 inst_15453 ( .A(net_9911), .Z(net_15301) );
NAND2_X2 inst_4205 ( .ZN(net_5290), .A1(net_5173), .A2(net_4979) );
CLKBUF_X2 inst_11452 ( .A(net_11299), .Z(net_11300) );
CLKBUF_X2 inst_9633 ( .A(net_9480), .Z(net_9481) );
CLKBUF_X2 inst_17039 ( .A(net_16886), .Z(net_16887) );
CLKBUF_X2 inst_17465 ( .A(net_17312), .Z(net_17313) );
CLKBUF_X2 inst_18747 ( .A(net_9231), .Z(net_18595) );
CLKBUF_X2 inst_12027 ( .A(net_9992), .Z(net_11875) );
CLKBUF_X2 inst_18265 ( .A(net_16984), .Z(net_18113) );
CLKBUF_X2 inst_18495 ( .A(net_18342), .Z(net_18343) );
CLKBUF_X2 inst_11063 ( .A(net_10910), .Z(net_10911) );
CLKBUF_X2 inst_9408 ( .A(net_9255), .Z(net_9256) );
INV_X4 inst_6156 ( .A(net_6198), .ZN(net_6197) );
CLKBUF_X2 inst_17999 ( .A(net_17846), .Z(net_17847) );
OAI21_X2 inst_3019 ( .B2(net_5044), .ZN(net_5041), .A(net_4886), .B1(net_1765) );
SDFFR_X2 inst_2327 ( .SE(net_2260), .Q(net_355), .D(net_355), .CK(net_11509), .RN(x6501), .SI(x2100) );
CLKBUF_X2 inst_13430 ( .A(net_13195), .Z(net_13278) );
INV_X4 inst_5078 ( .ZN(net_5846), .A(net_5791) );
DFFS_X2 inst_6866 ( .QN(net_6334), .D(net_5468), .CK(net_18932), .SN(x6501) );
CLKBUF_X2 inst_14976 ( .A(net_10333), .Z(net_14824) );
CLKBUF_X2 inst_11579 ( .A(net_11290), .Z(net_11427) );
XNOR2_X2 inst_113 ( .ZN(net_3925), .A(net_3543), .B(net_3542) );
CLKBUF_X2 inst_17212 ( .A(net_17059), .Z(net_17060) );
CLKBUF_X2 inst_10433 ( .A(net_10280), .Z(net_10281) );
CLKBUF_X2 inst_17217 ( .A(net_10461), .Z(net_17065) );
CLKBUF_X2 inst_16751 ( .A(net_15981), .Z(net_16599) );
CLKBUF_X2 inst_14023 ( .A(net_13870), .Z(net_13871) );
CLKBUF_X2 inst_9680 ( .A(net_9527), .Z(net_9528) );
AND2_X4 inst_9106 ( .ZN(net_2314), .A2(net_2082), .A1(net_2081) );
AOI22_X2 inst_8479 ( .B1(net_6609), .A1(net_6576), .A2(net_6257), .B2(net_6110), .ZN(net_3461) );
CLKBUF_X2 inst_10849 ( .A(net_10696), .Z(net_10697) );
CLKBUF_X2 inst_18633 ( .A(net_18480), .Z(net_18481) );
DFFR_X2 inst_7298 ( .QN(net_6325), .D(net_1142), .CK(net_14479), .RN(x6501) );
NAND2_X2 inst_4063 ( .ZN(net_5878), .A2(net_5765), .A1(net_3496) );
CLKBUF_X2 inst_10069 ( .A(net_9599), .Z(net_9917) );
AOI22_X2 inst_8340 ( .B1(net_8737), .A1(net_8515), .B2(net_4350), .A2(net_4349), .ZN(net_3707) );
CLKBUF_X2 inst_16427 ( .A(net_16274), .Z(net_16275) );
AOI211_X2 inst_9016 ( .C1(net_7303), .ZN(net_2022), .A(net_2021), .B(net_2020), .C2(net_2019) );
SDFFR_X2 inst_2625 ( .Q(net_7385), .D(net_7385), .SE(net_1136), .CK(net_18298), .RN(x6501), .SI(x4635) );
CLKBUF_X2 inst_14088 ( .A(net_13935), .Z(net_13936) );
INV_X4 inst_6064 ( .A(net_8295), .ZN(net_976) );
CLKBUF_X2 inst_19156 ( .A(net_19003), .Z(net_19004) );
CLKBUF_X2 inst_16081 ( .A(net_11592), .Z(net_15929) );
CLKBUF_X2 inst_12652 ( .A(net_12499), .Z(net_12500) );
CLKBUF_X2 inst_9244 ( .A(net_9091), .Z(net_9092) );
NOR2_X4 inst_3329 ( .ZN(net_3304), .A1(net_3159), .A2(net_3073) );
INV_X4 inst_5769 ( .A(net_7622), .ZN(net_557) );
CLKBUF_X2 inst_13844 ( .A(net_13691), .Z(net_13692) );
OR2_X4 inst_2847 ( .ZN(net_4316), .A1(net_1633), .A2(net_1632) );
SDFF_X2 inst_1442 ( .SI(net_7288), .Q(net_7105), .D(net_7105), .SE(net_6278), .CK(net_17713) );
XNOR2_X2 inst_332 ( .B(net_7639), .A(net_7636), .ZN(net_808) );
CLKBUF_X2 inst_14192 ( .A(net_14039), .Z(net_14040) );
NAND2_X4 inst_4013 ( .ZN(net_4642), .A1(net_4557), .A2(net_4506) );
SDFFR_X2 inst_2132 ( .SI(net_7199), .Q(net_7199), .D(net_6450), .SE(net_4362), .CK(net_14565), .RN(x6501) );
SDFF_X2 inst_1289 ( .Q(net_7828), .D(net_7828), .SE(net_2730), .SI(net_2712), .CK(net_17151) );
MUX2_X2 inst_4979 ( .A(net_9034), .Z(net_3974), .B(net_3269), .S(net_622) );
NAND2_X2 inst_4686 ( .A1(net_7166), .A2(net_2282), .ZN(net_2192) );
NAND2_X2 inst_4869 ( .ZN(net_1395), .A2(net_828), .A1(net_166) );
SDFF_X2 inst_1951 ( .D(net_7279), .SI(net_6936), .Q(net_6936), .SE(net_6281), .CK(net_18984) );
SDFF_X2 inst_378 ( .SI(net_8406), .Q(net_8406), .SE(net_3969), .D(net_3949), .CK(net_11026) );
CLKBUF_X2 inst_17831 ( .A(net_14005), .Z(net_17679) );
DFFR_X1 inst_7444 ( .QN(net_8924), .D(net_4759), .CK(net_14593), .RN(x6501) );
AOI22_X2 inst_8151 ( .B1(net_7916), .A1(net_7814), .B2(net_6103), .A2(net_4398), .ZN(net_4001) );
CLKBUF_X2 inst_11302 ( .A(net_11149), .Z(net_11150) );
CLKBUF_X2 inst_18205 ( .A(net_18052), .Z(net_18053) );
AOI221_X2 inst_8750 ( .B2(net_5657), .C2(net_5609), .ZN(net_5607), .A(net_5515), .B1(net_2699), .C1(net_366) );
SDFFR_X2 inst_2200 ( .SI(net_6484), .Q(net_6481), .D(net_6481), .SE(net_2897), .CK(net_9109), .RN(x6501) );
MUX2_X2 inst_4937 ( .Z(net_2853), .S(net_2852), .B(net_1918), .A(net_895) );
CLKBUF_X2 inst_10320 ( .A(net_10167), .Z(net_10168) );
AOI22_X2 inst_8284 ( .B1(net_8693), .A1(net_8656), .ZN(net_6228), .B2(net_6109), .A2(net_3857) );
AOI22_X2 inst_8080 ( .B1(net_8114), .A1(net_7876), .A2(net_6098), .B2(net_4190), .ZN(net_4065) );
CLKBUF_X2 inst_9948 ( .A(net_9795), .Z(net_9796) );
CLKBUF_X2 inst_14707 ( .A(net_14554), .Z(net_14555) );
XNOR2_X2 inst_250 ( .A(net_2729), .B(net_2681), .ZN(net_1200) );
CLKBUF_X2 inst_9275 ( .A(net_9077), .Z(net_9123) );
INV_X4 inst_5762 ( .A(net_6399), .ZN(net_1055) );
INV_X2 inst_6595 ( .A(net_6128), .ZN(net_6127) );
CLKBUF_X2 inst_9384 ( .A(net_9104), .Z(net_9232) );
SDFF_X2 inst_1523 ( .Q(net_7875), .D(net_7875), .SI(net_2585), .SE(net_2543), .CK(net_15841) );
CLKBUF_X2 inst_9941 ( .A(net_9788), .Z(net_9789) );
CLKBUF_X2 inst_17787 ( .A(net_17634), .Z(net_17635) );
SDFF_X2 inst_1048 ( .SI(net_7322), .Q(net_6696), .D(net_6696), .SE(net_3125), .CK(net_9158) );
DFFR_X2 inst_7120 ( .QN(net_7608), .D(net_3088), .CK(net_9797), .RN(x6501) );
CLKBUF_X2 inst_16822 ( .A(net_15969), .Z(net_16670) );
CLKBUF_X2 inst_18429 ( .A(net_12507), .Z(net_18277) );
CLKBUF_X2 inst_13537 ( .A(net_13384), .Z(net_13385) );
SDFFR_X2 inst_2270 ( .SI(net_7380), .SE(net_2793), .Q(net_239), .D(net_239), .CK(net_17832), .RN(x6501) );
CLKBUF_X2 inst_16050 ( .A(net_11551), .Z(net_15898) );
CLKBUF_X2 inst_11624 ( .A(net_11471), .Z(net_11472) );
SDFFR_X2 inst_2401 ( .SI(net_7371), .SE(net_2732), .D(net_2696), .QN(net_146), .CK(net_16107), .RN(x6501) );
CLKBUF_X2 inst_12979 ( .A(net_12826), .Z(net_12827) );
CLKBUF_X2 inst_10092 ( .A(net_9312), .Z(net_9940) );
CLKBUF_X2 inst_14723 ( .A(net_13501), .Z(net_14571) );
CLKBUF_X2 inst_12649 ( .A(net_12496), .Z(net_12497) );
CLKBUF_X2 inst_9356 ( .A(net_9203), .Z(net_9204) );
AOI22_X2 inst_8367 ( .B1(net_8888), .A1(net_8333), .B2(net_6252), .A2(net_4345), .ZN(net_3681) );
AOI22_X2 inst_8015 ( .B1(net_8167), .A1(net_7725), .B2(net_6101), .A2(net_6095), .ZN(net_6014) );
CLKBUF_X2 inst_15564 ( .A(net_15411), .Z(net_15412) );
AOI22_X2 inst_8196 ( .B1(net_8570), .A1(net_8459), .A2(net_6263), .B2(net_6262), .ZN(net_3840) );
INV_X4 inst_6050 ( .A(net_7360), .ZN(net_1284) );
CLKBUF_X2 inst_14287 ( .A(net_14134), .Z(net_14135) );
INV_X2 inst_6204 ( .ZN(net_5506), .A(net_5413) );
CLKBUF_X2 inst_17351 ( .A(net_12504), .Z(net_17199) );
AOI222_X1 inst_8618 ( .A2(net_8222), .ZN(net_4892), .A1(net_4891), .B1(net_4890), .B2(net_4889), .C2(net_4888), .C1(net_3133) );
CLKBUF_X2 inst_9710 ( .A(net_9122), .Z(net_9558) );
SDFF_X2 inst_420 ( .SI(net_8302), .Q(net_8302), .SE(net_3978), .D(net_3965), .CK(net_11113) );
NAND3_X2 inst_3992 ( .A2(net_8965), .A3(net_8901), .ZN(net_5036), .A1(net_1098) );
CLKBUF_X2 inst_12522 ( .A(net_12369), .Z(net_12370) );
NOR3_X2 inst_3265 ( .ZN(net_2842), .A1(net_2841), .A2(net_2840), .A3(net_2518) );
CLKBUF_X2 inst_15669 ( .A(net_14476), .Z(net_15517) );
DFFR_X1 inst_7558 ( .Q(net_7171), .D(net_6421), .CK(net_11845), .RN(x6501) );
SDFF_X2 inst_1305 ( .Q(net_7822), .D(net_7822), .SE(net_2730), .SI(net_2575), .CK(net_16082) );
AOI22_X2 inst_7997 ( .B1(net_8131), .A1(net_7893), .A2(net_6098), .B2(net_4190), .ZN(net_4136) );
XNOR2_X2 inst_314 ( .A(net_6829), .B(net_990), .ZN(net_951) );
CLKBUF_X2 inst_14813 ( .A(net_14660), .Z(net_14661) );
AOI221_X4 inst_8713 ( .C1(net_7938), .B1(net_7836), .C2(net_6103), .ZN(net_6049), .B2(net_4398), .A(net_4287) );
NOR4_X2 inst_3225 ( .ZN(net_2351), .A1(net_2111), .A2(net_1840), .A3(net_1491), .A4(net_1014) );
CLKBUF_X2 inst_13367 ( .A(net_12337), .Z(net_13215) );
CLKBUF_X2 inst_15342 ( .A(net_15189), .Z(net_15190) );
SDFF_X2 inst_597 ( .SI(net_8390), .Q(net_8390), .D(net_3974), .SE(net_3969), .CK(net_10836) );
INV_X4 inst_6161 ( .A(net_6251), .ZN(net_6250) );
INV_X4 inst_5524 ( .ZN(net_1356), .A(net_667) );
DFFR_X2 inst_7257 ( .QN(net_7404), .D(net_1975), .CK(net_17780), .RN(x6501) );
CLKBUF_X2 inst_11859 ( .A(net_10917), .Z(net_11707) );
DFFS_X1 inst_6927 ( .D(net_6145), .CK(net_16367), .SN(x6501), .Q(x845) );
CLKBUF_X2 inst_15115 ( .A(net_14962), .Z(net_14963) );
CLKBUF_X2 inst_12272 ( .A(net_12119), .Z(net_12120) );
CLKBUF_X2 inst_16985 ( .A(net_16832), .Z(net_16833) );
SDFF_X2 inst_472 ( .SI(net_8478), .Q(net_8478), .SE(net_3983), .D(net_3976), .CK(net_12799) );
SDFF_X2 inst_447 ( .Q(net_8777), .D(net_8777), .SE(net_3982), .SI(net_3948), .CK(net_13431) );
NAND2_X2 inst_4533 ( .ZN(net_3379), .A1(net_3378), .A2(net_3374) );
INV_X4 inst_5987 ( .A(net_8969), .ZN(net_1515) );
CLKBUF_X2 inst_12872 ( .A(net_10076), .Z(net_12720) );
CLKBUF_X2 inst_16940 ( .A(net_16787), .Z(net_16788) );
SDFFR_X2 inst_2623 ( .Q(net_7391), .D(net_2796), .SE(net_1136), .CK(net_18307), .RN(x6501), .SI(x4514) );
SDFF_X2 inst_1391 ( .SI(net_7714), .Q(net_7714), .D(net_2584), .SE(net_2559), .CK(net_16067) );
SDFF_X2 inst_665 ( .Q(net_8439), .D(net_8439), .SI(net_3951), .SE(net_3934), .CK(net_13409) );
NAND2_X2 inst_4843 ( .ZN(net_912), .A1(net_911), .A2(net_585) );
CLKBUF_X2 inst_16831 ( .A(net_16678), .Z(net_16679) );
CLKBUF_X2 inst_12929 ( .A(net_12776), .Z(net_12777) );
CLKBUF_X2 inst_12014 ( .A(net_9915), .Z(net_11862) );
CLKBUF_X2 inst_10219 ( .A(net_10066), .Z(net_10067) );
NOR2_X2 inst_3538 ( .A2(net_3162), .ZN(net_2643), .A1(net_811) );
NAND4_X2 inst_3755 ( .ZN(net_4266), .A1(net_3862), .A2(net_3859), .A3(net_3858), .A4(net_3856) );
AOI221_X4 inst_8718 ( .B1(net_8716), .C1(net_8494), .ZN(net_4351), .B2(net_4350), .C2(net_4349), .A(net_4264) );
CLKBUF_X2 inst_9810 ( .A(net_9657), .Z(net_9658) );
SDFF_X2 inst_1196 ( .SI(net_7300), .Q(net_7117), .D(net_7117), .SE(net_6278), .CK(net_18225) );
CLKBUF_X2 inst_17899 ( .A(net_13671), .Z(net_17747) );
CLKBUF_X2 inst_13815 ( .A(net_13662), .Z(net_13663) );
CLKBUF_X2 inst_18154 ( .A(net_16026), .Z(net_18002) );
NOR2_X2 inst_3428 ( .A2(net_3093), .ZN(net_3084), .A1(net_1186) );
CLKBUF_X2 inst_10510 ( .A(net_9656), .Z(net_10358) );
NOR2_X4 inst_3336 ( .A1(net_6106), .ZN(net_2327), .A2(net_2185) );
AOI22_X2 inst_7963 ( .B1(net_8092), .A1(net_7752), .B2(net_6108), .A2(net_6096), .ZN(net_4165) );
CLKBUF_X2 inst_19043 ( .A(net_17738), .Z(net_18891) );
AND4_X2 inst_9034 ( .ZN(net_5519), .A2(net_5023), .A4(net_4869), .A1(net_4780), .A3(net_4578) );
CLKBUF_X2 inst_16625 ( .A(net_16472), .Z(net_16473) );
OR2_X4 inst_2837 ( .ZN(net_2407), .A1(net_2406), .A2(net_2405) );
DFFR_X2 inst_7115 ( .QN(net_7609), .D(net_3055), .CK(net_9808), .RN(x6501) );
SDFF_X2 inst_1845 ( .D(net_7298), .SI(net_6915), .Q(net_6915), .SE(net_6284), .CK(net_18186) );
CLKBUF_X2 inst_17847 ( .A(net_17694), .Z(net_17695) );
CLKBUF_X2 inst_14681 ( .A(net_14528), .Z(net_14529) );
CLKBUF_X2 inst_9296 ( .A(net_9117), .Z(net_9144) );
CLKBUF_X2 inst_15598 ( .A(net_14145), .Z(net_15446) );
DFFS_X2 inst_6905 ( .QN(net_7525), .D(net_1798), .CK(net_16280), .SN(x6501) );
SDFF_X2 inst_1429 ( .SI(net_7265), .Q(net_7042), .D(net_7042), .SE(net_6280), .CK(net_17083) );
AOI22_X2 inst_8439 ( .B1(net_6600), .A1(net_6567), .A2(net_6257), .B2(net_6110), .ZN(net_3502) );
CLKBUF_X2 inst_12919 ( .A(net_11101), .Z(net_12767) );
SDFF_X2 inst_586 ( .Q(net_8821), .D(net_8821), .SE(net_3964), .SI(net_3947), .CK(net_12983) );
INV_X4 inst_5220 ( .ZN(net_2757), .A(net_2220) );
CLKBUF_X2 inst_9828 ( .A(net_9289), .Z(net_9676) );
DFFR_X2 inst_7176 ( .QN(net_7348), .D(net_2846), .CK(net_9563), .RN(x6501) );
CLKBUF_X2 inst_10563 ( .A(net_10410), .Z(net_10411) );
SDFFR_X2 inst_2591 ( .QN(net_7241), .D(net_2785), .SI(net_1945), .SE(net_1379), .CK(net_14744), .RN(x6501) );
CLKBUF_X2 inst_15317 ( .A(net_14466), .Z(net_15165) );
SDFFR_X1 inst_2652 ( .D(net_6756), .SE(net_4506), .CK(net_9331), .RN(x6501), .SI(x2195), .Q(x2195) );
INV_X4 inst_5221 ( .ZN(net_2685), .A(net_2220) );
SDFF_X2 inst_1203 ( .D(net_7300), .SI(net_6957), .Q(net_6957), .SE(net_6281), .CK(net_15916) );
SDFF_X2 inst_802 ( .SI(net_8341), .Q(net_8341), .D(net_3981), .SE(net_3880), .CK(net_10699) );
XNOR2_X2 inst_296 ( .B(net_7370), .ZN(net_986), .A(net_512) );
CLKBUF_X2 inst_16229 ( .A(net_16076), .Z(net_16077) );
CLKBUF_X2 inst_14626 ( .A(net_9339), .Z(net_14474) );
NAND2_X2 inst_4370 ( .A1(net_7073), .A2(net_5162), .ZN(net_5087) );
CLKBUF_X2 inst_11218 ( .A(net_11065), .Z(net_11066) );
AND2_X2 inst_9185 ( .ZN(net_2138), .A1(net_1930), .A2(net_1929) );
CLKBUF_X2 inst_11047 ( .A(net_10894), .Z(net_10895) );
NAND3_X2 inst_3943 ( .ZN(net_4471), .A1(net_4469), .A3(net_4468), .A2(net_4274) );
CLKBUF_X2 inst_14280 ( .A(net_14127), .Z(net_14128) );
SDFFR_X2 inst_2532 ( .SE(net_7164), .Q(net_7164), .D(net_2282), .SI(net_2146), .CK(net_18697), .RN(x6501) );
CLKBUF_X2 inst_13263 ( .A(net_13110), .Z(net_13111) );
SDFFR_X2 inst_2463 ( .QN(net_7413), .SE(net_3354), .SI(net_1468), .CK(net_10090), .D(x13984), .RN(x6501) );
CLKBUF_X2 inst_17267 ( .A(net_17114), .Z(net_17115) );
CLKBUF_X2 inst_11206 ( .A(net_11053), .Z(net_11054) );
CLKBUF_X2 inst_10907 ( .A(net_10754), .Z(net_10755) );
INV_X4 inst_5610 ( .A(net_7428), .ZN(net_3009) );
SDFF_X2 inst_1464 ( .SI(net_7301), .Q(net_7078), .D(net_7078), .SE(net_6280), .CK(net_15897) );
CLKBUF_X2 inst_15536 ( .A(net_12558), .Z(net_15384) );
CLKBUF_X2 inst_12778 ( .A(net_12625), .Z(net_12626) );
AOI22_X2 inst_8490 ( .B1(net_6678), .A1(net_6645), .A2(net_6213), .B2(net_6138), .ZN(net_3450) );
INV_X8 inst_5031 ( .ZN(net_5871), .A(net_5718) );
CLKBUF_X2 inst_19002 ( .A(net_18849), .Z(net_18850) );
CLKBUF_X2 inst_17656 ( .A(net_17503), .Z(net_17504) );
CLKBUF_X2 inst_13498 ( .A(net_13345), .Z(net_13346) );
CLKBUF_X2 inst_13215 ( .A(net_13062), .Z(net_13063) );
INV_X2 inst_6441 ( .ZN(net_624), .A(net_623) );
SDFF_X2 inst_1308 ( .SI(net_7700), .Q(net_7700), .SE(net_2714), .D(net_2704), .CK(net_14293) );
OAI21_X2 inst_3070 ( .B2(net_6456), .B1(net_4362), .ZN(net_4311), .A(net_2954) );
XOR2_X1 inst_85 ( .Z(net_2506), .A(net_2502), .B(net_1280) );
NAND2_X2 inst_4733 ( .ZN(net_2706), .A2(net_1586), .A1(net_1117) );
CLKBUF_X2 inst_16949 ( .A(net_16286), .Z(net_16797) );
INV_X4 inst_5963 ( .A(net_5976), .ZN(x3524) );
CLKBUF_X2 inst_14693 ( .A(net_14540), .Z(net_14541) );
CLKBUF_X2 inst_9681 ( .A(net_9353), .Z(net_9529) );
CLKBUF_X2 inst_16310 ( .A(net_16157), .Z(net_16158) );
CLKBUF_X2 inst_11850 ( .A(net_11697), .Z(net_11698) );
CLKBUF_X2 inst_12598 ( .A(net_12445), .Z(net_12446) );
CLKBUF_X2 inst_11314 ( .A(net_11161), .Z(net_11162) );
NAND2_X4 inst_4022 ( .A1(net_3573), .ZN(net_3562), .A2(net_3561) );
SDFF_X2 inst_1978 ( .D(net_7280), .SI(net_7017), .Q(net_7017), .SE(net_6277), .CK(net_18978) );
XNOR2_X2 inst_290 ( .B(net_7380), .ZN(net_1002), .A(net_525) );
CLKBUF_X2 inst_15285 ( .A(net_15132), .Z(net_15133) );
CLKBUF_X2 inst_16346 ( .A(net_13838), .Z(net_16194) );
CLKBUF_X2 inst_14122 ( .A(net_13969), .Z(net_13970) );
SDFFR_X2 inst_2112 ( .SE(net_5582), .D(net_5523), .CK(net_14206), .RN(x6501), .SI(x52), .Q(x52) );
AOI22_X2 inst_7743 ( .B1(net_6972), .A1(net_6932), .A2(net_5443), .B2(net_5442), .ZN(net_5434) );
CLKBUF_X2 inst_16610 ( .A(net_16457), .Z(net_16458) );
CLKBUF_X2 inst_15431 ( .A(net_15278), .Z(net_15279) );
OAI21_X2 inst_3036 ( .B2(net_8231), .B1(net_4928), .ZN(net_4842), .A(net_3545) );
SDFF_X2 inst_814 ( .SI(net_8504), .Q(net_8504), .D(net_3963), .SE(net_3884), .CK(net_10897) );
CLKBUF_X2 inst_13441 ( .A(net_13288), .Z(net_13289) );
CLKBUF_X2 inst_9465 ( .A(net_9312), .Z(net_9313) );
CLKBUF_X2 inst_19007 ( .A(net_13394), .Z(net_18855) );
INV_X4 inst_5203 ( .ZN(net_2428), .A(net_2427) );
AOI21_X2 inst_8973 ( .ZN(net_2468), .A(net_2467), .B2(net_2466), .B1(net_791) );
NOR2_X2 inst_3471 ( .ZN(net_2438), .A2(net_2280), .A1(net_1736) );
SDFF_X2 inst_1458 ( .SI(net_7278), .Q(net_7135), .D(net_7135), .SE(net_6279), .CK(net_14637) );
CLKBUF_X2 inst_15933 ( .A(net_12262), .Z(net_15781) );
CLKBUF_X2 inst_11332 ( .A(net_11179), .Z(net_11180) );
SDFFR_X2 inst_2275 ( .SI(net_7387), .SE(net_2814), .Q(net_246), .D(net_246), .CK(net_14714), .RN(x6501) );
CLKBUF_X2 inst_16650 ( .A(net_10676), .Z(net_16498) );
CLKBUF_X2 inst_15727 ( .A(net_15574), .Z(net_15575) );
CLKBUF_X2 inst_10212 ( .A(net_10059), .Z(net_10060) );
CLKBUF_X2 inst_16567 ( .A(net_11748), .Z(net_16415) );
SDFF_X2 inst_822 ( .SI(net_8514), .Q(net_8514), .D(net_3950), .SE(net_3884), .CK(net_10513) );
CLKBUF_X2 inst_12053 ( .A(net_11011), .Z(net_11901) );
SDFF_X2 inst_1125 ( .D(net_7312), .SI(net_6554), .Q(net_6554), .SE(net_3070), .CK(net_11998) );
NAND2_X2 inst_4341 ( .A1(net_7145), .A2(net_5166), .ZN(net_5116) );
INV_X4 inst_5996 ( .A(net_7662), .ZN(net_1645) );
CLKBUF_X2 inst_10984 ( .A(net_10831), .Z(net_10832) );
SDFF_X2 inst_609 ( .SI(net_8404), .Q(net_8404), .D(net_3976), .SE(net_3969), .CK(net_12539) );
CLKBUF_X2 inst_11521 ( .A(net_11136), .Z(net_11369) );
AOI22_X2 inst_8261 ( .B1(net_8689), .A1(net_8652), .B2(net_6109), .A2(net_3857), .ZN(net_3777) );
SDFF_X2 inst_795 ( .SI(net_8367), .Q(net_8367), .D(net_3976), .SE(net_3880), .CK(net_12515) );
SDFFR_X2 inst_2491 ( .Q(net_8985), .D(net_8985), .SI(net_2626), .SE(net_2562), .CK(net_14533), .RN(x6501) );
HA_X1 inst_6668 ( .S(net_3229), .CO(net_3228), .A(net_3227), .B(net_3090) );
CLKBUF_X2 inst_14127 ( .A(net_13974), .Z(net_13975) );
CLKBUF_X2 inst_11179 ( .A(net_10186), .Z(net_11027) );
CLKBUF_X2 inst_12848 ( .A(net_12571), .Z(net_12696) );
AOI22_X2 inst_8215 ( .B1(net_8868), .A1(net_8313), .B2(net_6252), .A2(net_4345), .ZN(net_3821) );
SDFF_X2 inst_619 ( .SI(net_8530), .Q(net_8530), .SE(net_3979), .D(net_3962), .CK(net_13117) );
CLKBUF_X2 inst_14481 ( .A(net_14328), .Z(net_14329) );
CLKBUF_X2 inst_12139 ( .A(net_11986), .Z(net_11987) );
SDFF_X2 inst_1654 ( .SI(net_7707), .Q(net_7707), .D(net_2655), .SE(net_2559), .CK(net_15504) );
NAND2_X2 inst_4547 ( .A1(net_3378), .ZN(net_3317), .A2(net_3315) );
AOI22_X2 inst_7831 ( .A2(net_5535), .B2(net_5260), .ZN(net_4690), .B1(net_3056), .A1(net_455) );
CLKBUF_X2 inst_10545 ( .A(net_10235), .Z(net_10393) );
CLKBUF_X2 inst_10553 ( .A(net_10400), .Z(net_10401) );
CLKBUF_X2 inst_10265 ( .A(net_10112), .Z(net_10113) );
INV_X2 inst_6486 ( .A(net_9051), .ZN(net_904) );
SDFFS_X2 inst_2076 ( .SE(net_2794), .SI(net_2785), .Q(net_170), .D(net_170), .CK(net_14938), .SN(x6501) );
CLKBUF_X2 inst_18896 ( .A(net_18743), .Z(net_18744) );
INV_X4 inst_5879 ( .A(net_7423), .ZN(net_3014) );
CLKBUF_X2 inst_16835 ( .A(net_16682), .Z(net_16683) );
SDFFR_X2 inst_2481 ( .Q(net_8991), .D(net_8991), .SI(net_2606), .SE(net_2562), .CK(net_17270), .RN(x6501) );
AOI22_X2 inst_7824 ( .A2(net_5535), .B2(net_5260), .ZN(net_4700), .B1(net_4699), .A1(net_447) );
CLKBUF_X2 inst_11474 ( .A(net_9694), .Z(net_11322) );
CLKBUF_X2 inst_13385 ( .A(net_13232), .Z(net_13233) );
NAND2_X2 inst_4285 ( .A1(net_6887), .A2(net_5247), .ZN(net_5175) );
CLKBUF_X2 inst_15386 ( .A(net_9737), .Z(net_15234) );
SDFF_X2 inst_1162 ( .SI(net_7316), .Q(net_6591), .D(net_6591), .SE(net_3069), .CK(net_12070) );
CLKBUF_X2 inst_18829 ( .A(net_18676), .Z(net_18677) );
DFFR_X1 inst_7485 ( .QN(net_7426), .D(net_4042), .CK(net_12377), .RN(x6501) );
CLKBUF_X2 inst_14384 ( .A(net_14231), .Z(net_14232) );
INV_X4 inst_6108 ( .ZN(net_2700), .A(net_155) );
INV_X2 inst_6572 ( .ZN(net_828), .A(net_210) );
CLKBUF_X2 inst_13123 ( .A(net_12970), .Z(net_12971) );
DFFR_X1 inst_7449 ( .QN(net_8932), .D(net_4750), .CK(net_17313), .RN(x6501) );
OAI221_X2 inst_2973 ( .C2(net_2489), .B2(net_2450), .ZN(net_2419), .A(net_2273), .C1(net_1271), .B1(net_736) );
CLKBUF_X2 inst_11454 ( .A(net_11301), .Z(net_11302) );
CLKBUF_X2 inst_17297 ( .A(net_12197), .Z(net_17145) );
SDFF_X2 inst_1433 ( .SI(net_7263), .Q(net_7080), .D(net_7080), .SE(net_6278), .CK(net_14368) );
SDFF_X2 inst_793 ( .SI(net_8364), .Q(net_8364), .D(net_3940), .SE(net_3880), .CK(net_10236) );
CLKBUF_X2 inst_18923 ( .A(net_18770), .Z(net_18771) );
NAND2_X2 inst_4815 ( .ZN(net_1249), .A2(net_902), .A1(net_782) );
SDFF_X2 inst_1999 ( .SI(net_7911), .Q(net_7911), .D(net_2655), .SE(net_2461), .CK(net_15383) );
SDFFR_X1 inst_2733 ( .SI(net_9046), .Q(net_9046), .D(net_7475), .SE(net_3208), .CK(net_12208), .RN(x6501) );
CLKBUF_X2 inst_12405 ( .A(net_11408), .Z(net_12253) );
CLKBUF_X2 inst_11750 ( .A(net_11597), .Z(net_11598) );
CLKBUF_X2 inst_15429 ( .A(net_15276), .Z(net_15277) );
AOI221_X2 inst_8808 ( .C2(net_5535), .B2(net_5260), .A(net_4898), .ZN(net_4720), .B1(net_661), .C1(net_473) );
CLKBUF_X2 inst_17225 ( .A(net_9643), .Z(net_17073) );
SDFF_X2 inst_475 ( .SI(net_8448), .Q(net_8448), .SE(net_3983), .D(net_3977), .CK(net_12471) );
CLKBUF_X2 inst_13253 ( .A(net_12488), .Z(net_13101) );
CLKBUF_X2 inst_9436 ( .A(net_9283), .Z(net_9284) );
CLKBUF_X2 inst_19020 ( .A(net_18867), .Z(net_18868) );
CLKBUF_X2 inst_17958 ( .A(net_17805), .Z(net_17806) );
NAND2_X2 inst_4738 ( .ZN(net_2749), .A2(net_1586), .A1(net_1033) );
CLKBUF_X2 inst_9412 ( .A(net_9222), .Z(net_9260) );
CLKBUF_X2 inst_17917 ( .A(net_12608), .Z(net_17765) );
NAND2_X2 inst_4412 ( .A1(net_6851), .A2(net_5016), .ZN(net_5015) );
CLKBUF_X2 inst_12595 ( .A(net_10772), .Z(net_12443) );
CLKBUF_X2 inst_9564 ( .A(net_9411), .Z(net_9412) );
CLKBUF_X2 inst_12804 ( .A(net_12651), .Z(net_12652) );
CLKBUF_X2 inst_15573 ( .A(net_15420), .Z(net_15421) );
INV_X4 inst_5724 ( .A(net_7261), .ZN(net_567) );
AOI22_X2 inst_8276 ( .A1(net_8617), .B1(net_8432), .A2(net_3864), .B2(net_3863), .ZN(net_3765) );
NAND2_X2 inst_4331 ( .A1(net_7061), .A2(net_5162), .ZN(net_5126) );
CLKBUF_X2 inst_11054 ( .A(net_10458), .Z(net_10902) );
AOI22_X2 inst_8049 ( .B1(net_8205), .A1(net_7695), .B2(net_6099), .A2(net_4399), .ZN(net_4091) );
NAND2_X2 inst_4705 ( .ZN(net_2713), .A2(net_1586), .A1(net_927) );
CLKBUF_X2 inst_10940 ( .A(net_9513), .Z(net_10788) );
CLKBUF_X2 inst_11543 ( .A(net_10577), .Z(net_11391) );
CLKBUF_X2 inst_16178 ( .A(net_16025), .Z(net_16026) );
CLKBUF_X2 inst_16320 ( .A(net_12274), .Z(net_16168) );
NOR2_X2 inst_3580 ( .A2(net_7625), .ZN(net_1077), .A1(net_565) );
CLKBUF_X2 inst_12321 ( .A(net_12168), .Z(net_12169) );
CLKBUF_X2 inst_11531 ( .A(net_9469), .Z(net_11379) );
CLKBUF_X2 inst_10004 ( .A(net_9851), .Z(net_9852) );
OAI21_X2 inst_3080 ( .ZN(net_3256), .A(net_3186), .B2(net_3185), .B1(net_3080) );
DFF_X1 inst_6857 ( .Q(net_6426), .D(net_3624), .CK(net_17954) );
CLKBUF_X2 inst_19181 ( .A(net_19028), .Z(net_19029) );
SDFFR_X2 inst_2434 ( .D(net_4890), .SE(net_2683), .SI(net_405), .Q(net_405), .CK(net_13834), .RN(x6501) );
DFFR_X1 inst_7432 ( .QN(net_8912), .D(net_4855), .CK(net_16694), .RN(x6501) );
SDFF_X2 inst_1107 ( .D(net_7338), .SI(net_6547), .Q(net_6547), .SE(net_3086), .CK(net_9464) );
CLKBUF_X2 inst_10039 ( .A(net_9469), .Z(net_9887) );
CLKBUF_X2 inst_15335 ( .A(net_14550), .Z(net_15183) );
CLKBUF_X2 inst_12909 ( .A(net_10683), .Z(net_12757) );
INV_X4 inst_5930 ( .A(net_8291), .ZN(net_999) );
CLKBUF_X2 inst_9916 ( .A(net_9491), .Z(net_9764) );
CLKBUF_X2 inst_18288 ( .A(net_18135), .Z(net_18136) );
NAND2_X2 inst_4253 ( .A1(net_6909), .A2(net_5247), .ZN(net_5207) );
SDFFR_X1 inst_2776 ( .D(net_7396), .Q(net_7293), .SI(net_1939), .SE(net_1327), .CK(net_15374), .RN(x6501) );
CLKBUF_X2 inst_9646 ( .A(net_9493), .Z(net_9494) );
AOI222_X1 inst_8612 ( .B2(net_6758), .B1(net_5835), .A2(net_5830), .C2(net_5824), .ZN(net_5801), .C1(net_2130), .A1(net_1219) );
SDFF_X2 inst_746 ( .Q(net_8794), .D(net_8794), .SI(net_3944), .SE(net_3879), .CK(net_12260) );
CLKBUF_X2 inst_13016 ( .A(net_12863), .Z(net_12864) );
INV_X2 inst_6553 ( .A(net_7214), .ZN(net_501) );
CLKBUF_X2 inst_17618 ( .A(net_17465), .Z(net_17466) );
AOI222_X1 inst_8660 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3906), .B1(net_3271), .C1(net_3269), .A1(x13750) );
SDFFR_X2 inst_2267 ( .SI(net_7377), .SE(net_2793), .Q(net_236), .D(net_236), .CK(net_13711), .RN(x6501) );
CLKBUF_X2 inst_18722 ( .A(net_18569), .Z(net_18570) );
DFFR_X2 inst_7127 ( .QN(net_7604), .D(net_3075), .CK(net_9786), .RN(x6501) );
CLKBUF_X2 inst_18019 ( .A(net_14081), .Z(net_17867) );
CLKBUF_X2 inst_17664 ( .A(net_17511), .Z(net_17512) );
INV_X4 inst_5662 ( .A(net_7368), .ZN(net_936) );
AOI22_X2 inst_7893 ( .B1(net_9002), .A2(net_5538), .B2(net_5456), .ZN(net_4536), .A1(net_431) );
CLKBUF_X2 inst_16299 ( .A(net_12119), .Z(net_16147) );
CLKBUF_X2 inst_10050 ( .A(net_9897), .Z(net_9898) );
INV_X4 inst_5820 ( .A(net_7610), .ZN(net_2829) );
AOI221_X4 inst_8721 ( .B1(net_8721), .C1(net_8499), .B2(net_4350), .C2(net_4349), .ZN(net_4346), .A(net_4259) );
SDFF_X2 inst_1577 ( .Q(net_8029), .D(net_8029), .SI(net_2722), .SE(net_2545), .CK(net_18384) );
SDFF_X2 inst_1110 ( .D(net_7341), .SI(net_6550), .Q(net_6550), .SE(net_3086), .CK(net_11871) );
INV_X4 inst_5778 ( .A(net_9057), .ZN(net_622) );
CLKBUF_X2 inst_18607 ( .A(net_18454), .Z(net_18455) );
CLKBUF_X2 inst_14870 ( .A(net_14717), .Z(net_14718) );
OR2_X2 inst_2873 ( .ZN(net_4511), .A1(net_4510), .A2(net_4509) );
AOI22_X2 inst_8468 ( .B1(net_6540), .A1(net_6507), .A2(net_6137), .B2(net_6104), .ZN(net_3472) );
SDFFR_X2 inst_2442 ( .D(net_2669), .SE(net_2313), .SI(net_407), .Q(net_407), .CK(net_16530), .RN(x6501) );
CLKBUF_X2 inst_9676 ( .A(net_9523), .Z(net_9524) );
SDFFS_X2 inst_2066 ( .SI(net_7392), .SE(net_2417), .Q(net_181), .D(net_181), .CK(net_17744), .SN(x6501) );
CLKBUF_X2 inst_12126 ( .A(net_11973), .Z(net_11974) );
SDFF_X2 inst_1742 ( .Q(net_8137), .D(net_8137), .SI(net_2711), .SE(net_2541), .CK(net_16986) );
CLKBUF_X2 inst_12085 ( .A(net_11932), .Z(net_11933) );
CLKBUF_X2 inst_13603 ( .A(net_13450), .Z(net_13451) );
CLKBUF_X2 inst_12091 ( .A(net_10776), .Z(net_11939) );
CLKBUF_X2 inst_18282 ( .A(net_14824), .Z(net_18130) );
INV_X2 inst_6236 ( .ZN(net_5454), .A(net_5273) );
CLKBUF_X2 inst_18843 ( .A(net_17938), .Z(net_18691) );
CLKBUF_X2 inst_18903 ( .A(net_18750), .Z(net_18751) );
NAND2_X2 inst_4779 ( .ZN(net_1613), .A1(net_1612), .A2(net_1327) );
CLKBUF_X2 inst_9522 ( .A(net_9221), .Z(net_9370) );
CLKBUF_X2 inst_19010 ( .A(net_18857), .Z(net_18858) );
OAI211_X4 inst_3175 ( .ZN(net_5987), .C2(net_5985), .C1(net_5984), .B(net_2514), .A(net_2169) );
SDFFR_X2 inst_2302 ( .D(net_2750), .SE(net_2683), .SI(net_465), .Q(net_465), .CK(net_16926), .RN(x6501) );
CLKBUF_X2 inst_11021 ( .A(net_10868), .Z(net_10869) );
CLKBUF_X2 inst_16289 ( .A(net_16136), .Z(net_16137) );
CLKBUF_X2 inst_9967 ( .A(net_9228), .Z(net_9815) );
DFFR_X2 inst_7181 ( .QN(net_8952), .D(net_2468), .CK(net_17235), .RN(x6501) );
SDFFR_X2 inst_2447 ( .D(net_3309), .SE(net_2313), .SI(net_413), .Q(net_413), .CK(net_13932), .RN(x6501) );
CLKBUF_X2 inst_12043 ( .A(net_11890), .Z(net_11891) );
CLKBUF_X2 inst_17377 ( .A(net_15168), .Z(net_17225) );
CLKBUF_X2 inst_18393 ( .A(net_18240), .Z(net_18241) );
CLKBUF_X2 inst_11648 ( .A(net_9891), .Z(net_11496) );
CLKBUF_X2 inst_15408 ( .A(net_15255), .Z(net_15256) );
CLKBUF_X2 inst_11151 ( .A(net_9834), .Z(net_10999) );
CLKBUF_X2 inst_10914 ( .A(net_10761), .Z(net_10762) );
CLKBUF_X2 inst_9695 ( .A(net_9212), .Z(net_9543) );
INV_X4 inst_6141 ( .A(net_6121), .ZN(net_6120) );
AOI22_X2 inst_7921 ( .A1(net_8989), .A2(net_5456), .B2(net_5260), .ZN(net_4461), .B1(net_3272) );
CLKBUF_X2 inst_13303 ( .A(net_13150), .Z(net_13151) );
DFFR_X2 inst_7163 ( .QN(net_6396), .D(net_2756), .CK(net_18949), .RN(x6501) );
NAND2_X2 inst_4803 ( .A2(net_2255), .ZN(net_1500), .A1(net_757) );
SDFF_X2 inst_935 ( .SI(net_7342), .Q(net_6683), .D(net_6683), .SE(net_3126), .CK(net_11690) );
CLKBUF_X2 inst_17860 ( .A(net_17707), .Z(net_17708) );
INV_X2 inst_6619 ( .A(net_6251), .ZN(net_6249) );
INV_X4 inst_5699 ( .A(net_7414), .ZN(net_1039) );
NAND2_X2 inst_4772 ( .A1(net_6324), .A2(net_2307), .ZN(net_2075) );
CLKBUF_X2 inst_12781 ( .A(net_12628), .Z(net_12629) );
NAND2_X2 inst_4634 ( .ZN(net_2646), .A2(net_2480), .A1(net_2479) );
CLKBUF_X2 inst_16655 ( .A(net_15851), .Z(net_16503) );
CLKBUF_X2 inst_11255 ( .A(net_9903), .Z(net_11103) );
CLKBUF_X2 inst_15997 ( .A(net_15844), .Z(net_15845) );
CLKBUF_X2 inst_9284 ( .A(net_9131), .Z(net_9132) );
CLKBUF_X2 inst_11587 ( .A(net_11434), .Z(net_11435) );
OAI22_X2 inst_2944 ( .A1(net_2043), .ZN(net_1798), .A2(net_1797), .B2(net_1136), .B1(net_685) );
INV_X8 inst_5011 ( .ZN(net_5657), .A(net_4413) );
CLKBUF_X2 inst_15830 ( .A(net_15677), .Z(net_15678) );
CLKBUF_X2 inst_15186 ( .A(net_9361), .Z(net_15034) );
CLKBUF_X2 inst_13690 ( .A(net_13537), .Z(net_13538) );
CLKBUF_X2 inst_18972 ( .A(net_9896), .Z(net_18820) );
AOI22_X2 inst_8314 ( .A1(net_8595), .B1(net_8410), .A2(net_3864), .B2(net_3863), .ZN(net_3731) );
OR2_X4 inst_2862 ( .ZN(net_6283), .A2(net_2199), .A1(net_805) );
AOI22_X2 inst_7949 ( .B1(net_7920), .A1(net_7818), .B2(net_6103), .A2(net_4398), .ZN(net_4177) );
AOI22_X2 inst_8391 ( .B1(net_8673), .A1(net_8636), .B2(net_6109), .A2(net_3857), .ZN(net_3658) );
CLKBUF_X2 inst_13397 ( .A(net_9384), .Z(net_13245) );
CLKBUF_X2 inst_15109 ( .A(net_11465), .Z(net_14957) );
INV_X2 inst_6510 ( .ZN(net_534), .A(x13271) );
INV_X4 inst_5808 ( .A(net_8962), .ZN(net_2309) );
CLKBUF_X2 inst_16132 ( .A(net_14897), .Z(net_15980) );
CLKBUF_X2 inst_12181 ( .A(net_12028), .Z(net_12029) );
CLKBUF_X2 inst_13390 ( .A(net_9298), .Z(net_13238) );
CLKBUF_X2 inst_11268 ( .A(net_10767), .Z(net_11116) );
DFFS_X2 inst_6859 ( .Q(net_6321), .D(net_5524), .CK(net_17464), .SN(x6501) );
DFFR_X1 inst_7439 ( .Q(net_7516), .D(net_4843), .CK(net_13606), .RN(x6501) );
NAND2_X2 inst_4454 ( .A2(net_4962), .ZN(net_4961), .A1(net_3253) );
CLKBUF_X2 inst_17342 ( .A(net_16873), .Z(net_17190) );
CLKBUF_X2 inst_12813 ( .A(net_12660), .Z(net_12661) );
AOI221_X4 inst_8709 ( .C1(net_7934), .B1(net_7832), .C2(net_6103), .ZN(net_6041), .B2(net_4398), .A(net_4292) );
NAND2_X2 inst_4315 ( .A1(net_7097), .A2(net_5164), .ZN(net_5142) );
SDFF_X2 inst_365 ( .SI(net_8522), .Q(net_8522), .SE(net_3979), .D(net_3977), .CK(net_11117) );
XOR2_X1 inst_67 ( .Z(net_4208), .A(net_3579), .B(x2451) );
SDFF_X2 inst_954 ( .SI(net_7313), .Q(net_6687), .D(net_6687), .SE(net_3125), .CK(net_12046) );
CLKBUF_X2 inst_16436 ( .A(net_16283), .Z(net_16284) );
CLKBUF_X2 inst_13162 ( .A(net_13009), .Z(net_13010) );
CLKBUF_X2 inst_16844 ( .A(net_16691), .Z(net_16692) );
CLKBUF_X2 inst_14186 ( .A(net_14033), .Z(net_14034) );
CLKBUF_X2 inst_11216 ( .A(net_11063), .Z(net_11064) );
AOI22_X2 inst_8569 ( .A2(net_8250), .A1(net_4729), .B2(net_4728), .B1(net_2790), .ZN(net_2155) );
CLKBUF_X2 inst_17729 ( .A(net_17576), .Z(net_17577) );
CLKBUF_X2 inst_11685 ( .A(net_11532), .Z(net_11533) );
SDFF_X2 inst_1823 ( .D(net_7263), .SI(net_6840), .Q(net_6840), .SE(net_6282), .CK(net_14349) );
INV_X4 inst_5084 ( .ZN(net_5730), .A(net_5709) );
XNOR2_X2 inst_202 ( .ZN(net_1541), .B(net_1200), .A(net_1185) );
CLKBUF_X2 inst_16249 ( .A(net_16096), .Z(net_16097) );
DFFR_X2 inst_7359 ( .Q(net_7330), .CK(net_9532), .D(x13011), .RN(x6501) );
AND2_X2 inst_9154 ( .ZN(net_2972), .A2(net_2971), .A1(net_1154) );
SDFFR_X2 inst_2212 ( .Q(net_7445), .D(net_7445), .SE(net_2863), .CK(net_12820), .SI(x13619), .RN(x6501) );
CLKBUF_X2 inst_13786 ( .A(net_10975), .Z(net_13634) );
SDFF_X2 inst_1401 ( .Q(net_8191), .D(net_8191), .SI(net_2706), .SE(net_2561), .CK(net_18059) );
NAND2_X2 inst_4830 ( .ZN(net_1318), .A2(net_1078), .A1(net_572) );
CLKBUF_X2 inst_13444 ( .A(net_12781), .Z(net_13292) );
SDFF_X2 inst_2030 ( .SI(net_7924), .Q(net_7924), .D(net_2575), .SE(net_2461), .CK(net_16014) );
AOI22_X2 inst_8254 ( .B1(net_8836), .A1(net_8355), .A2(net_6265), .B2(net_6253), .ZN(net_6064) );
CLKBUF_X2 inst_11172 ( .A(net_11019), .Z(net_11020) );
XOR2_X2 inst_30 ( .A(net_6796), .Z(net_1210), .B(net_1209) );
SDFF_X2 inst_610 ( .SI(net_8405), .Q(net_8405), .SE(net_3969), .D(net_3939), .CK(net_10543) );
INV_X2 inst_6271 ( .A(net_4553), .ZN(net_4509) );
CLKBUF_X2 inst_16107 ( .A(net_12590), .Z(net_15955) );
XNOR2_X2 inst_233 ( .ZN(net_1251), .B(net_865), .A(net_495) );
CLKBUF_X2 inst_9704 ( .A(net_9102), .Z(net_9552) );
AOI222_X1 inst_8639 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3985), .B1(net_2820), .C1(net_2818), .A1(x13833) );
AOI222_X1 inst_8595 ( .B2(net_6772), .B1(net_5835), .ZN(net_5833), .C2(net_5832), .A2(net_5830), .A1(net_3104), .C1(x2948) );
CLKBUF_X2 inst_17852 ( .A(net_17699), .Z(net_17700) );
CLKBUF_X2 inst_12296 ( .A(net_12143), .Z(net_12144) );
CLKBUF_X2 inst_9527 ( .A(net_9286), .Z(net_9375) );
AND2_X4 inst_9127 ( .A1(net_2742), .ZN(net_1295), .A2(x14005) );
CLKBUF_X2 inst_18822 ( .A(net_18669), .Z(net_18670) );
XOR2_X2 inst_60 ( .A(net_3224), .Z(net_952), .B(net_588) );
AOI21_X2 inst_8939 ( .B2(net_5871), .ZN(net_5660), .A(net_5659), .B1(net_2688) );
INV_X16 inst_6651 ( .ZN(net_6261), .A(net_4456) );
CLKBUF_X2 inst_13540 ( .A(net_11783), .Z(net_13388) );
AOI22_X2 inst_7752 ( .B1(net_6980), .A1(net_6940), .A2(net_5443), .B2(net_5442), .ZN(net_5398) );
CLKBUF_X2 inst_13285 ( .A(net_13132), .Z(net_13133) );
CLKBUF_X2 inst_12862 ( .A(net_12709), .Z(net_12710) );
DFFR_X2 inst_7339 ( .Q(net_7327), .CK(net_11772), .D(x13031), .RN(x6501) );
CLKBUF_X2 inst_12189 ( .A(net_12036), .Z(net_12037) );
CLKBUF_X2 inst_10392 ( .A(net_10239), .Z(net_10240) );
AOI22_X2 inst_8389 ( .B1(net_8784), .A1(net_8525), .ZN(net_6234), .A2(net_3861), .B2(net_3860) );
CLKBUF_X2 inst_14397 ( .A(net_14244), .Z(net_14245) );
NOR2_X2 inst_3478 ( .ZN(net_2406), .A2(net_2245), .A1(net_834) );
CLKBUF_X2 inst_18727 ( .A(net_18574), .Z(net_18575) );
CLKBUF_X2 inst_11252 ( .A(net_11099), .Z(net_11100) );
CLKBUF_X2 inst_10181 ( .A(net_9542), .Z(net_10029) );
CLKBUF_X2 inst_17238 ( .A(net_17085), .Z(net_17086) );
DFFR_X2 inst_7147 ( .QN(net_7167), .D(net_3035), .CK(net_15206), .RN(x6501) );
CLKBUF_X2 inst_15505 ( .A(net_14475), .Z(net_15353) );
SDFFR_X1 inst_2782 ( .D(net_7383), .Q(net_7280), .SI(net_1961), .SE(net_1327), .CK(net_18160), .RN(x6501) );
DFFR_X2 inst_7248 ( .QN(net_7258), .D(net_2051), .CK(net_15187), .RN(x6501) );
INV_X4 inst_5475 ( .A(net_1716), .ZN(net_872) );
CLKBUF_X2 inst_13887 ( .A(net_13734), .Z(net_13735) );
CLKBUF_X2 inst_11191 ( .A(net_11038), .Z(net_11039) );
NAND4_X2 inst_3720 ( .ZN(net_4310), .A1(net_4197), .A2(net_4196), .A3(net_4195), .A4(net_4194) );
CLKBUF_X2 inst_14672 ( .A(net_10361), .Z(net_14520) );
CLKBUF_X2 inst_11964 ( .A(net_11039), .Z(net_11812) );
CLKBUF_X2 inst_12444 ( .A(net_9089), .Z(net_12292) );
SDFF_X2 inst_2005 ( .SI(net_7782), .Q(net_7782), .D(net_2584), .SE(net_2459), .CK(net_16016) );
CLKBUF_X2 inst_11988 ( .A(net_11835), .Z(net_11836) );
CLKBUF_X2 inst_13377 ( .A(net_12738), .Z(net_13225) );
SDFF_X2 inst_736 ( .SI(net_8355), .Q(net_8355), .D(net_3956), .SE(net_3880), .CK(net_13238) );
SDFF_X2 inst_544 ( .Q(net_8687), .D(net_8687), .SI(net_3957), .SE(net_3935), .CK(net_11016) );
INV_X4 inst_5865 ( .A(net_8926), .ZN(net_2608) );
AOI22_X2 inst_8021 ( .B1(net_8201), .A1(net_7691), .B2(net_6099), .A2(net_4399), .ZN(net_4115) );
INV_X4 inst_5465 ( .ZN(net_760), .A(net_759) );
AOI22_X2 inst_8232 ( .A1(net_8612), .B1(net_8427), .A2(net_3864), .B2(net_3863), .ZN(net_3805) );
CLKBUF_X2 inst_17290 ( .A(net_17137), .Z(net_17138) );
NAND2_X2 inst_4402 ( .A1(net_7087), .A2(net_5164), .ZN(net_5055) );
SDFF_X2 inst_734 ( .SI(net_8363), .Q(net_8363), .D(net_3952), .SE(net_3880), .CK(net_10339) );
DFFR_X2 inst_7352 ( .Q(net_7328), .CK(net_11768), .D(x13025), .RN(x6501) );
SDFF_X2 inst_1282 ( .Q(net_7831), .D(net_7831), .SE(net_2730), .SI(net_2711), .CK(net_17096) );
AOI22_X2 inst_8528 ( .B1(net_6524), .A1(net_6491), .A2(net_6137), .B2(net_6104), .ZN(net_3412) );
CLKBUF_X2 inst_16125 ( .A(net_15972), .Z(net_15973) );
CLKBUF_X2 inst_14818 ( .A(net_14665), .Z(net_14666) );
CLKBUF_X2 inst_15673 ( .A(net_15520), .Z(net_15521) );
CLKBUF_X2 inst_17715 ( .A(net_12266), .Z(net_17563) );
CLKBUF_X2 inst_10425 ( .A(net_10075), .Z(net_10273) );
AOI21_X2 inst_8898 ( .ZN(net_5865), .A(net_5783), .B1(net_5662), .B2(net_5037) );
CLKBUF_X2 inst_19033 ( .A(net_18880), .Z(net_18881) );
INV_X4 inst_5634 ( .A(net_7563), .ZN(net_2936) );
CLKBUF_X2 inst_9597 ( .A(net_9444), .Z(net_9445) );
NOR2_X2 inst_3587 ( .A1(net_6793), .ZN(net_6170), .A2(net_1897) );
AOI221_X2 inst_8777 ( .B2(net_5657), .C2(net_5535), .ZN(net_5262), .A(net_4918), .B1(net_2733), .C1(net_445) );
CLKBUF_X2 inst_10139 ( .A(net_9986), .Z(net_9987) );
CLKBUF_X2 inst_13003 ( .A(net_12850), .Z(net_12851) );
CLKBUF_X2 inst_10147 ( .A(net_9994), .Z(net_9995) );
CLKBUF_X2 inst_18053 ( .A(net_17900), .Z(net_17901) );
INV_X4 inst_5543 ( .ZN(net_645), .A(x3079) );
INV_X2 inst_6392 ( .A(net_7630), .ZN(net_1181) );
CLKBUF_X2 inst_17706 ( .A(net_17553), .Z(net_17554) );
INV_X4 inst_5588 ( .A(net_7380), .ZN(net_1462) );
CLKBUF_X2 inst_15465 ( .A(net_15312), .Z(net_15313) );
CLKBUF_X2 inst_11427 ( .A(net_11274), .Z(net_11275) );
CLKBUF_X2 inst_16203 ( .A(net_16050), .Z(net_16051) );
INV_X2 inst_6183 ( .ZN(net_5841), .A(net_5786) );
CLKBUF_X2 inst_17800 ( .A(net_17647), .Z(net_17648) );
CLKBUF_X2 inst_11529 ( .A(net_11376), .Z(net_11377) );
AOI22_X2 inst_8542 ( .B1(net_6660), .A1(net_6627), .A2(net_6213), .B2(net_6138), .ZN(net_3398) );
CLKBUF_X2 inst_17745 ( .A(net_17592), .Z(net_17593) );
CLKBUF_X2 inst_16445 ( .A(net_16292), .Z(net_16293) );
NAND4_X2 inst_3701 ( .A4(net_6228), .A1(net_6227), .ZN(net_4436), .A2(net_3757), .A3(net_3756) );
NOR2_X2 inst_3357 ( .ZN(net_5568), .A1(net_5400), .A2(net_5399) );
DFFR_X2 inst_7082 ( .QN(net_7662), .D(net_3895), .CK(net_12681), .RN(x6501) );
CLKBUF_X2 inst_11822 ( .A(net_11669), .Z(net_11670) );
XOR2_X2 inst_8 ( .Z(net_2498), .B(net_2494), .A(net_2464) );
CLKBUF_X2 inst_15559 ( .A(net_15406), .Z(net_15407) );
CLKBUF_X2 inst_15456 ( .A(net_14184), .Z(net_15304) );
AOI21_X2 inst_8925 ( .A(net_5745), .ZN(net_5721), .B2(net_5584), .B1(net_4872) );
DFFR_X2 inst_6984 ( .QN(net_5958), .D(net_5895), .CK(net_9230), .RN(x6501) );
CLKBUF_X2 inst_17420 ( .A(net_17267), .Z(net_17268) );
SDFFS_X2 inst_2090 ( .D(net_6835), .SI(net_6829), .Q(net_6829), .SE(net_2146), .CK(net_18677), .SN(x6501) );
SDFF_X2 inst_965 ( .SI(net_7324), .Q(net_6731), .D(net_6731), .SE(net_3124), .CK(net_9884) );
AOI22_X2 inst_8228 ( .B1(net_8833), .A1(net_8352), .A2(net_6265), .B2(net_6253), .ZN(net_3809) );
CLKBUF_X2 inst_14583 ( .A(net_14430), .Z(net_14431) );
CLKBUF_X2 inst_12267 ( .A(net_12114), .Z(net_12115) );
AOI222_X1 inst_8677 ( .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3310), .C1(net_3309), .B1(net_3143), .A2(net_3106) );
CLKBUF_X2 inst_11991 ( .A(net_11838), .Z(net_11839) );
CLKBUF_X2 inst_12284 ( .A(net_12131), .Z(net_12132) );
CLKBUF_X2 inst_11976 ( .A(net_10359), .Z(net_11824) );
INV_X4 inst_5392 ( .ZN(net_1317), .A(net_1082) );
INV_X2 inst_6179 ( .ZN(net_5885), .A(net_5884) );
CLKBUF_X2 inst_15520 ( .A(net_11722), .Z(net_15368) );
CLKBUF_X2 inst_18073 ( .A(net_17920), .Z(net_17921) );
CLKBUF_X2 inst_16003 ( .A(net_15850), .Z(net_15851) );
AOI22_X2 inst_7913 ( .B1(net_8972), .B2(net_5456), .A2(net_4501), .ZN(net_4500), .A1(net_2742) );
CLKBUF_X2 inst_16097 ( .A(net_15944), .Z(net_15945) );
CLKBUF_X2 inst_13288 ( .A(net_13135), .Z(net_13136) );
CLKBUF_X2 inst_14013 ( .A(net_13860), .Z(net_13861) );
SDFF_X2 inst_1934 ( .SI(net_8045), .Q(net_8045), .D(net_2585), .SE(net_2508), .CK(net_15732) );
DFF_X1 inst_6759 ( .Q(net_7538), .D(net_4614), .CK(net_11977) );
CLKBUF_X2 inst_16022 ( .A(net_12509), .Z(net_15870) );
CLKBUF_X2 inst_9429 ( .A(net_9113), .Z(net_9277) );
CLKBUF_X2 inst_18207 ( .A(net_9799), .Z(net_18055) );
NAND3_X2 inst_3916 ( .ZN(net_5622), .A1(net_5551), .A3(net_5485), .A2(net_5328) );
INV_X4 inst_5739 ( .A(net_7347), .ZN(net_1085) );
INV_X4 inst_5401 ( .ZN(net_1113), .A(net_881) );
CLKBUF_X2 inst_18752 ( .A(net_18599), .Z(net_18600) );
CLKBUF_X2 inst_9970 ( .A(net_9817), .Z(net_9818) );
CLKBUF_X2 inst_17007 ( .A(net_16854), .Z(net_16855) );
AOI22_X2 inst_8319 ( .B1(net_8697), .A1(net_8660), .ZN(net_6232), .B2(net_6109), .A2(net_3857) );
AOI22_X2 inst_8539 ( .B1(net_6593), .A1(net_6560), .A2(net_6257), .B2(net_6110), .ZN(net_3401) );
CLKBUF_X2 inst_19136 ( .A(net_18983), .Z(net_18984) );
CLKBUF_X2 inst_13359 ( .A(net_13206), .Z(net_13207) );
AOI22_X2 inst_8464 ( .B1(net_6587), .A1(net_6554), .A2(net_6257), .B2(net_6110), .ZN(net_3476) );
CLKBUF_X2 inst_10968 ( .A(net_10815), .Z(net_10816) );
SDFFS_X2 inst_2097 ( .Q(net_7524), .D(net_7524), .SI(net_4956), .SE(net_1136), .CK(net_18902), .SN(x6501) );
CLKBUF_X2 inst_12943 ( .A(net_12790), .Z(net_12791) );
NAND2_X2 inst_4484 ( .A2(net_5267), .ZN(net_4494), .A1(net_169) );
CLKBUF_X2 inst_14948 ( .A(net_14795), .Z(net_14796) );
AOI22_X2 inst_8053 ( .B1(net_8070), .A1(net_7866), .B2(net_6107), .A2(net_4400), .ZN(net_4088) );
INV_X2 inst_6215 ( .ZN(net_5495), .A(net_5369) );
CLKBUF_X2 inst_18798 ( .A(net_18645), .Z(net_18646) );
CLKBUF_X2 inst_16350 ( .A(net_14554), .Z(net_16198) );
CLKBUF_X2 inst_16700 ( .A(net_10739), .Z(net_16548) );
CLKBUF_X2 inst_12225 ( .A(net_12072), .Z(net_12073) );
SDFF_X2 inst_1050 ( .SI(net_7339), .Q(net_6680), .D(net_6680), .SE(net_3126), .CK(net_11891) );
INV_X2 inst_6476 ( .ZN(net_920), .A(net_221) );
CLKBUF_X2 inst_17546 ( .A(net_17393), .Z(net_17394) );
CLKBUF_X2 inst_17195 ( .A(net_16541), .Z(net_17043) );
NAND2_X2 inst_4661 ( .ZN(net_2464), .A1(net_2232), .A2(net_2231) );
SDFF_X2 inst_1852 ( .D(net_7275), .SI(net_6932), .Q(net_6932), .SE(net_6281), .CK(net_17357) );
DFF_X1 inst_6809 ( .Q(net_8226), .D(net_4419), .CK(net_17224) );
INV_X2 inst_6273 ( .ZN(net_4378), .A(net_4366) );
NOR3_X2 inst_3282 ( .ZN(net_2386), .A1(net_2385), .A3(net_2318), .A2(net_1877) );
CLKBUF_X2 inst_12667 ( .A(net_12514), .Z(net_12515) );
NAND2_X2 inst_4074 ( .A2(net_6766), .A1(net_5835), .ZN(net_5772) );
NAND4_X2 inst_3783 ( .ZN(net_4238), .A1(net_3684), .A2(net_3683), .A3(net_3682), .A4(net_3681) );
CLKBUF_X2 inst_13613 ( .A(net_9970), .Z(net_13461) );
SDFF_X2 inst_1557 ( .Q(net_8022), .D(net_8022), .SI(net_2574), .SE(net_2545), .CK(net_15589) );
SDFFR_X2 inst_2399 ( .SI(net_7368), .SE(net_2732), .D(net_2698), .QN(net_143), .CK(net_16115), .RN(x6501) );
CLKBUF_X2 inst_18498 ( .A(net_13699), .Z(net_18346) );
CLKBUF_X2 inst_18430 ( .A(net_18277), .Z(net_18278) );
CLKBUF_X2 inst_12207 ( .A(net_12054), .Z(net_12055) );
NOR2_X2 inst_3412 ( .A1(net_8896), .ZN(net_3325), .A2(net_3230) );
NAND2_X2 inst_4698 ( .A2(net_2315), .ZN(net_2223), .A1(net_1885) );
CLKBUF_X2 inst_9620 ( .A(net_9467), .Z(net_9468) );
AOI22_X2 inst_8485 ( .B1(net_6743), .A1(net_6710), .B2(net_6202), .A2(net_3520), .ZN(net_3455) );
CLKBUF_X2 inst_17431 ( .A(net_17278), .Z(net_17279) );
CLKBUF_X2 inst_17247 ( .A(net_17094), .Z(net_17095) );
CLKBUF_X2 inst_11326 ( .A(net_11173), .Z(net_11174) );
SDFF_X2 inst_1616 ( .Q(net_8157), .D(net_8157), .SI(net_2706), .SE(net_2538), .CK(net_18858) );
CLKBUF_X2 inst_14090 ( .A(net_13937), .Z(net_13938) );
AOI221_X2 inst_8813 ( .C2(net_5535), .A(net_5520), .B2(net_5260), .ZN(net_4715), .B1(net_4714), .C1(net_452) );
INV_X4 inst_5646 ( .A(net_8215), .ZN(net_742) );
CLKBUF_X2 inst_13167 ( .A(net_13014), .Z(net_13015) );
CLKBUF_X2 inst_11295 ( .A(net_10942), .Z(net_11143) );
CLKBUF_X2 inst_11403 ( .A(net_11250), .Z(net_11251) );
INV_X4 inst_5356 ( .ZN(net_1309), .A(net_1149) );
CLKBUF_X2 inst_13110 ( .A(net_12957), .Z(net_12958) );
AOI222_X1 inst_8690 ( .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3273), .C1(net_3272), .B1(net_3140), .A2(net_3109) );
CLKBUF_X2 inst_11786 ( .A(net_11633), .Z(net_11634) );
CLKBUF_X2 inst_11621 ( .A(net_11468), .Z(net_11469) );
CLKBUF_X2 inst_17410 ( .A(net_17257), .Z(net_17258) );
CLKBUF_X2 inst_15303 ( .A(net_15150), .Z(net_15151) );
CLKBUF_X2 inst_16536 ( .A(net_14401), .Z(net_16384) );
OAI211_X2 inst_3186 ( .ZN(net_5024), .B(net_4957), .A(net_4684), .C2(net_4554), .C1(net_1880) );
CLKBUF_X2 inst_15266 ( .A(net_15113), .Z(net_15114) );
NAND4_X2 inst_3762 ( .ZN(net_4259), .A1(net_3817), .A2(net_3816), .A3(net_3815), .A4(net_3814) );
INV_X4 inst_5653 ( .A(net_7394), .ZN(net_1864) );
CLKBUF_X2 inst_10925 ( .A(net_10772), .Z(net_10773) );
NOR3_X2 inst_3259 ( .A3(net_6209), .ZN(net_4397), .A2(net_1584), .A1(net_1380) );
SDFF_X2 inst_854 ( .SI(net_8634), .Q(net_8634), .D(net_3938), .SE(net_3885), .CK(net_12943) );
CLKBUF_X2 inst_12464 ( .A(net_10009), .Z(net_12312) );
CLKBUF_X2 inst_13293 ( .A(net_13140), .Z(net_13141) );
CLKBUF_X2 inst_13796 ( .A(net_13643), .Z(net_13644) );
CLKBUF_X2 inst_15369 ( .A(net_13583), .Z(net_15217) );
CLKBUF_X2 inst_16600 ( .A(net_16447), .Z(net_16448) );
NAND4_X2 inst_3678 ( .A4(net_6028), .A1(net_6027), .ZN(net_4587), .A2(net_4022), .A3(net_4021) );
NAND3_X2 inst_3979 ( .A1(net_6156), .ZN(net_2245), .A3(net_872), .A2(net_483) );
INV_X2 inst_6297 ( .ZN(net_4201), .A(net_3910) );
CLKBUF_X2 inst_15578 ( .A(net_15425), .Z(net_15426) );
AOI22_X2 inst_7865 ( .B2(net_5609), .A2(net_5267), .ZN(net_4576), .B1(net_380), .A1(net_184) );
CLKBUF_X2 inst_10478 ( .A(net_10325), .Z(net_10326) );
CLKBUF_X2 inst_12006 ( .A(net_11853), .Z(net_11854) );
AOI22_X2 inst_8008 ( .B1(net_8030), .A1(net_7996), .B2(net_6102), .A2(net_6097), .ZN(net_6040) );
CLKBUF_X2 inst_13401 ( .A(net_13248), .Z(net_13249) );
CLKBUF_X2 inst_10861 ( .A(net_9662), .Z(net_10709) );
CLKBUF_X2 inst_9464 ( .A(net_9311), .Z(net_9312) );
SDFF_X2 inst_1749 ( .SI(net_7289), .Q(net_7146), .D(net_7146), .SE(net_6279), .CK(net_15344) );
CLKBUF_X2 inst_16508 ( .A(net_16355), .Z(net_16356) );
CLKBUF_X2 inst_9717 ( .A(net_9564), .Z(net_9565) );
INV_X2 inst_6519 ( .ZN(net_804), .A(net_216) );
CLKBUF_X2 inst_14105 ( .A(net_12012), .Z(net_13953) );
INV_X4 inst_5514 ( .ZN(net_679), .A(net_678) );
CLKBUF_X2 inst_12518 ( .A(net_12365), .Z(net_12366) );
AND2_X4 inst_9071 ( .ZN(net_6257), .A2(net_3248), .A1(net_3216) );
CLKBUF_X2 inst_11872 ( .A(net_9253), .Z(net_11720) );
AOI211_X2 inst_9017 ( .ZN(net_2157), .A(net_1928), .C1(net_1927), .B(net_1649), .C2(net_892) );
SDFF_X2 inst_840 ( .SI(net_8650), .Q(net_8650), .D(net_3957), .SE(net_3885), .CK(net_10977) );
CLKBUF_X2 inst_16555 ( .A(net_16402), .Z(net_16403) );
CLKBUF_X2 inst_17073 ( .A(net_16920), .Z(net_16921) );
CLKBUF_X2 inst_11900 ( .A(net_11747), .Z(net_11748) );
CLKBUF_X2 inst_13523 ( .A(net_13370), .Z(net_13371) );
CLKBUF_X2 inst_12498 ( .A(net_11770), .Z(net_12346) );
INV_X4 inst_6117 ( .A(net_7404), .ZN(net_669) );
CLKBUF_X2 inst_10736 ( .A(net_10583), .Z(net_10584) );
INV_X4 inst_5876 ( .A(net_8917), .ZN(net_4736) );
DFFR_X1 inst_7497 ( .QN(net_6403), .D(net_3024), .CK(net_18017), .RN(x6501) );
NAND2_X2 inst_4294 ( .A1(net_7090), .ZN(net_5165), .A2(net_5164) );
CLKBUF_X2 inst_18512 ( .A(net_18359), .Z(net_18360) );
CLKBUF_X2 inst_14302 ( .A(net_14149), .Z(net_14150) );
CLKBUF_X2 inst_10799 ( .A(net_9662), .Z(net_10647) );
INV_X4 inst_5710 ( .A(net_6391), .ZN(net_1583) );
CLKBUF_X2 inst_9536 ( .A(net_9383), .Z(net_9384) );
INV_X4 inst_5939 ( .A(net_7253), .ZN(net_1960) );
CLKBUF_X2 inst_15966 ( .A(net_15813), .Z(net_15814) );
CLKBUF_X2 inst_11846 ( .A(net_11693), .Z(net_11694) );
INV_X4 inst_5679 ( .A(net_7651), .ZN(net_3595) );
DFFR_X2 inst_7272 ( .QN(net_7230), .D(net_1983), .CK(net_14775), .RN(x6501) );
CLKBUF_X2 inst_11141 ( .A(net_10988), .Z(net_10989) );
AND2_X2 inst_9200 ( .ZN(net_6085), .A2(net_1306), .A1(x13291) );
CLKBUF_X2 inst_16527 ( .A(net_16374), .Z(net_16375) );
SDFF_X2 inst_617 ( .SI(net_8519), .Q(net_8519), .SE(net_3979), .D(net_3961), .CK(net_13198) );
CLKBUF_X2 inst_14897 ( .A(net_9311), .Z(net_14745) );
AND2_X2 inst_9167 ( .ZN(net_2806), .A2(net_2553), .A1(net_1073) );
INV_X4 inst_5734 ( .A(net_7306), .ZN(net_1237) );
CLKBUF_X2 inst_10823 ( .A(net_10670), .Z(net_10671) );
CLKBUF_X2 inst_18089 ( .A(net_17936), .Z(net_17937) );
CLKBUF_X2 inst_16634 ( .A(net_16481), .Z(net_16482) );
AOI22_X2 inst_8123 ( .B1(net_7912), .A1(net_7810), .B2(net_6103), .A2(net_4398), .ZN(net_4026) );
INV_X2 inst_6614 ( .A(net_6206), .ZN(net_6205) );
CLKBUF_X2 inst_18457 ( .A(net_18304), .Z(net_18305) );
CLKBUF_X2 inst_15749 ( .A(net_15596), .Z(net_15597) );
INV_X4 inst_6029 ( .A(net_7391), .ZN(net_672) );
CLKBUF_X2 inst_19089 ( .A(net_18936), .Z(net_18937) );
CLKBUF_X2 inst_11956 ( .A(net_11803), .Z(net_11804) );
INV_X4 inst_5482 ( .A(net_1612), .ZN(net_734) );
DFFR_X2 inst_7159 ( .QN(net_5948), .D(net_2784), .CK(net_11220), .RN(x6501) );
DFF_X1 inst_6739 ( .Q(net_6784), .D(net_5630), .CK(net_9200) );
CLKBUF_X2 inst_17494 ( .A(net_17341), .Z(net_17342) );
CLKBUF_X2 inst_18045 ( .A(net_17892), .Z(net_17893) );
AOI21_X2 inst_8916 ( .ZN(net_5762), .A(net_5745), .B2(net_5596), .B1(net_4791) );
CLKBUF_X2 inst_14487 ( .A(net_14334), .Z(net_14335) );
CLKBUF_X2 inst_9818 ( .A(net_9665), .Z(net_9666) );
AOI221_X2 inst_8798 ( .C2(net_6187), .B2(net_5609), .A(net_4898), .ZN(net_4879), .B1(net_369), .C1(net_193) );
CLKBUF_X2 inst_15064 ( .A(net_14911), .Z(net_14912) );
OAI22_X2 inst_2909 ( .A2(net_8231), .B2(net_6133), .A1(net_4954), .ZN(net_4875), .B1(net_1411) );
CLKBUF_X2 inst_12636 ( .A(net_9762), .Z(net_12484) );
OAI21_X2 inst_3135 ( .ZN(net_2065), .B2(net_2060), .A(net_1970), .B1(net_641) );
SDFF_X2 inst_701 ( .Q(net_8429), .D(net_8429), .SI(net_3956), .SE(net_3934), .CK(net_13244) );
SDFFR_X2 inst_2380 ( .SE(net_2260), .Q(net_335), .D(net_335), .CK(net_9292), .RN(x6501), .SI(x2400) );
CLKBUF_X2 inst_16780 ( .A(net_16627), .Z(net_16628) );
CLKBUF_X2 inst_12337 ( .A(net_12184), .Z(net_12185) );
DFFR_X1 inst_7583 ( .Q(net_6827), .D(net_6815), .CK(net_15116), .RN(x6501) );
INV_X4 inst_5261 ( .ZN(net_2127), .A(net_1771) );
CLKBUF_X2 inst_15998 ( .A(net_15845), .Z(net_15846) );
CLKBUF_X2 inst_17356 ( .A(net_17203), .Z(net_17204) );
AOI22_X2 inst_7739 ( .A2(net_6755), .B2(net_6198), .ZN(net_5836), .A1(net_5835), .B1(x3651) );
DFFS_X1 inst_6933 ( .D(net_6145), .CK(net_16352), .SN(x6501), .Q(x879) );
SDFF_X2 inst_1007 ( .D(net_7319), .SI(net_6627), .Q(net_6627), .SE(net_3123), .CK(net_12029) );
CLKBUF_X2 inst_11011 ( .A(net_9120), .Z(net_10859) );
CLKBUF_X2 inst_15989 ( .A(net_13173), .Z(net_15837) );
CLKBUF_X2 inst_11674 ( .A(net_11521), .Z(net_11522) );
CLKBUF_X2 inst_11932 ( .A(net_11779), .Z(net_11780) );
INV_X4 inst_5066 ( .ZN(net_5910), .A(net_5864) );
CLKBUF_X2 inst_11998 ( .A(net_9293), .Z(net_11846) );
CLKBUF_X2 inst_16160 ( .A(net_16007), .Z(net_16008) );
OR2_X2 inst_2883 ( .ZN(net_1901), .A1(net_1900), .A2(net_1899) );
CLKBUF_X2 inst_11313 ( .A(net_10656), .Z(net_11161) );
CLKBUF_X2 inst_11108 ( .A(net_10955), .Z(net_10956) );
CLKBUF_X2 inst_18733 ( .A(net_14065), .Z(net_18581) );
CLKBUF_X2 inst_10083 ( .A(net_9930), .Z(net_9931) );
NAND4_X2 inst_3685 ( .A4(net_6244), .A1(net_6243), .ZN(net_4452), .A2(net_3855), .A3(net_3854) );
CLKBUF_X2 inst_10527 ( .A(net_10374), .Z(net_10375) );
CLKBUF_X2 inst_16407 ( .A(net_13049), .Z(net_16255) );
DFFS_X2 inst_6891 ( .QN(net_8968), .D(net_2857), .CK(net_17617), .SN(x6501) );
CLKBUF_X2 inst_11301 ( .A(net_11148), .Z(net_11149) );
CLKBUF_X2 inst_19140 ( .A(net_17292), .Z(net_18988) );
SDFF_X2 inst_1472 ( .SI(net_7302), .Q(net_7159), .D(net_7159), .SE(net_6279), .CK(net_15896) );
CLKBUF_X2 inst_19161 ( .A(net_17838), .Z(net_19009) );
CLKBUF_X2 inst_17633 ( .A(net_17480), .Z(net_17481) );
NAND2_X2 inst_4261 ( .A1(net_6912), .A2(net_5247), .ZN(net_5199) );
CLKBUF_X2 inst_12511 ( .A(net_12358), .Z(net_12359) );
CLKBUF_X2 inst_14784 ( .A(net_9880), .Z(net_14632) );
NAND4_X2 inst_3784 ( .ZN(net_4237), .A1(net_3677), .A2(net_3676), .A3(net_3675), .A4(net_3674) );
SDFF_X2 inst_1183 ( .SI(net_7327), .Q(net_6602), .D(net_6602), .SE(net_3069), .CK(net_9830) );
CLKBUF_X2 inst_9577 ( .A(net_9424), .Z(net_9425) );
SDFF_X2 inst_1489 ( .SI(net_7285), .Q(net_7102), .D(net_7102), .SE(net_6278), .CK(net_19025) );
SDFFR_X2 inst_2415 ( .D(net_2689), .SE(net_2313), .SI(net_459), .Q(net_459), .CK(net_13943), .RN(x6501) );
CLKBUF_X2 inst_12353 ( .A(net_12200), .Z(net_12201) );
CLKBUF_X2 inst_14498 ( .A(net_14345), .Z(net_14346) );
MUX2_X2 inst_4981 ( .A(net_9033), .Z(net_3958), .B(net_3098), .S(net_622) );
AOI22_X2 inst_8352 ( .B1(net_8849), .A1(net_8368), .A2(net_6265), .B2(net_6253), .ZN(net_3696) );
INV_X4 inst_5506 ( .ZN(net_2843), .A(net_692) );
DFFR_X2 inst_7102 ( .QN(net_5980), .D(net_3244), .CK(net_11229), .RN(x6501) );
SDFF_X2 inst_1808 ( .D(net_7291), .SI(net_6948), .Q(net_6948), .SE(net_6281), .CK(net_15338) );
CLKBUF_X2 inst_17896 ( .A(net_17743), .Z(net_17744) );
AOI22_X2 inst_8440 ( .B1(net_6534), .A1(net_6501), .A2(net_6137), .B2(net_6104), .ZN(net_3501) );
SDFF_X2 inst_988 ( .D(net_7325), .SI(net_6633), .Q(net_6633), .SE(net_3123), .CK(net_9165) );
CLKBUF_X2 inst_16988 ( .A(net_16835), .Z(net_16836) );
CLKBUF_X2 inst_10288 ( .A(net_9905), .Z(net_10136) );
CLKBUF_X2 inst_15668 ( .A(net_15515), .Z(net_15516) );
CLKBUF_X2 inst_14941 ( .A(net_14788), .Z(net_14789) );
CLKBUF_X2 inst_9333 ( .A(net_9180), .Z(net_9181) );
MUX2_X2 inst_4954 ( .A(net_2785), .S(net_2376), .Z(net_2369), .B(net_887) );
NAND2_X2 inst_4308 ( .A1(net_7135), .A2(net_5166), .ZN(net_5149) );
CLKBUF_X2 inst_11026 ( .A(net_10251), .Z(net_10874) );
CLKBUF_X2 inst_18460 ( .A(net_16965), .Z(net_18308) );
DFFR_X1 inst_7569 ( .Q(net_8287), .D(net_8277), .CK(net_11256), .RN(x6501) );
CLKBUF_X2 inst_18100 ( .A(net_17658), .Z(net_17948) );
CLKBUF_X2 inst_18654 ( .A(net_18501), .Z(net_18502) );
CLKBUF_X2 inst_10049 ( .A(net_9808), .Z(net_9897) );
CLKBUF_X2 inst_15249 ( .A(net_12077), .Z(net_15097) );
CLKBUF_X2 inst_9808 ( .A(net_9655), .Z(net_9656) );
INV_X4 inst_5527 ( .ZN(net_3233), .A(net_663) );
DFFR_X2 inst_7007 ( .QN(net_6309), .D(net_5798), .CK(net_16946), .RN(x6501) );
DFF_X1 inst_6718 ( .Q(net_6755), .D(net_5651), .CK(net_10448) );
CLKBUF_X2 inst_12562 ( .A(net_12231), .Z(net_12410) );
INV_X4 inst_5919 ( .ZN(net_2694), .A(net_160) );
CLKBUF_X2 inst_13471 ( .A(net_13318), .Z(net_13319) );
CLKBUF_X2 inst_17910 ( .A(net_17757), .Z(net_17758) );
CLKBUF_X2 inst_18939 ( .A(net_13260), .Z(net_18787) );
NAND2_X2 inst_4618 ( .A2(net_6144), .ZN(net_2605), .A1(net_2604) );
DFF_X1 inst_6827 ( .Q(net_6447), .D(net_3621), .CK(net_17917) );
SDFF_X2 inst_1922 ( .D(net_7268), .SI(net_6965), .Q(net_6965), .SE(net_6283), .CK(net_14325) );
NOR2_X2 inst_3361 ( .ZN(net_5564), .A1(net_5384), .A2(net_5383) );
OAI21_X2 inst_3170 ( .B2(net_2569), .ZN(net_1263), .B1(net_1262), .A(net_884) );
NOR4_X2 inst_3232 ( .A1(net_2309), .ZN(net_2076), .A3(net_2075), .A4(net_1869), .A2(net_1061) );
AOI22_X2 inst_8335 ( .B1(net_8810), .A1(net_8551), .A2(net_3861), .B2(net_3860), .ZN(net_3712) );
CLKBUF_X2 inst_13062 ( .A(net_12041), .Z(net_12910) );
CLKBUF_X2 inst_10524 ( .A(net_10371), .Z(net_10372) );
CLKBUF_X2 inst_10444 ( .A(net_10291), .Z(net_10292) );
INV_X4 inst_5973 ( .A(net_5964), .ZN(x3028) );
DFFS_X1 inst_6942 ( .D(net_6145), .CK(net_13640), .SN(x6501), .Q(x753) );
CLKBUF_X2 inst_16731 ( .A(net_16578), .Z(net_16579) );
SDFF_X2 inst_1350 ( .Q(net_8196), .D(net_8196), .SI(net_2575), .SE(net_2561), .CK(net_16002) );
CLKBUF_X2 inst_12156 ( .A(net_12003), .Z(net_12004) );
CLKBUF_X2 inst_16489 ( .A(net_16336), .Z(net_16337) );
OAI21_X2 inst_3012 ( .ZN(net_5740), .A(net_5718), .B2(net_5540), .B1(net_4975) );
CLKBUF_X2 inst_11369 ( .A(net_11216), .Z(net_11217) );
SDFFR_X2 inst_2635 ( .Q(net_7396), .D(net_7396), .SE(net_1136), .CK(net_15791), .RN(x6501), .SI(x4448) );
CLKBUF_X2 inst_16502 ( .A(net_16349), .Z(net_16350) );
CLKBUF_X2 inst_14014 ( .A(net_13861), .Z(net_13862) );
AOI222_X1 inst_8673 ( .C2(net_5832), .A2(net_5830), .B2(net_5824), .ZN(net_3496), .A1(net_3201), .B1(net_2041), .C1(x2261) );
NOR2_X2 inst_3363 ( .ZN(net_5562), .A1(net_5376), .A2(net_5375) );
SDFFR_X1 inst_2666 ( .D(net_6763), .SE(net_4506), .CK(net_9326), .RN(x6501), .SI(x1977), .Q(x1977) );
DFFR_X2 inst_7188 ( .QN(net_6420), .D(net_2432), .CK(net_18663), .RN(x6501) );
SDFF_X2 inst_1357 ( .SI(net_7752), .Q(net_7752), .D(net_2589), .SE(net_2560), .CK(net_18406) );
CLKBUF_X2 inst_18969 ( .A(net_18816), .Z(net_18817) );
CLKBUF_X2 inst_10938 ( .A(net_10785), .Z(net_10786) );
CLKBUF_X2 inst_9547 ( .A(net_9119), .Z(net_9395) );
INV_X4 inst_5302 ( .A(net_1704), .ZN(net_1689) );
NAND2_X2 inst_4476 ( .A2(net_5595), .ZN(net_4558), .A1(net_319) );
CLKBUF_X2 inst_11307 ( .A(net_11154), .Z(net_11155) );
DFFS_X2 inst_6861 ( .Q(net_6320), .D(net_5526), .CK(net_17463), .SN(x6501) );
SDFFR_X2 inst_2288 ( .SI(net_7482), .Q(net_7482), .D(net_2760), .SE(net_2441), .CK(net_16133), .RN(x6501) );
CLKBUF_X2 inst_13644 ( .A(net_12593), .Z(net_13492) );
CLKBUF_X2 inst_11505 ( .A(net_11352), .Z(net_11353) );
NAND2_X2 inst_4841 ( .A2(net_7358), .A1(net_1908), .ZN(net_1292) );
CLKBUF_X2 inst_9368 ( .A(net_9215), .Z(net_9216) );
SDFF_X2 inst_1834 ( .D(net_7267), .SI(net_6844), .Q(net_6844), .SE(net_6282), .CK(net_14118) );
CLKBUF_X2 inst_18870 ( .A(net_17335), .Z(net_18718) );
CLKBUF_X2 inst_17989 ( .A(net_17836), .Z(net_17837) );
NOR2_X2 inst_3574 ( .ZN(net_3326), .A2(net_1151), .A1(net_1075) );
SDFFR_X2 inst_2228 ( .Q(net_7472), .D(net_7472), .SE(net_2863), .CK(net_12176), .SI(x13414), .RN(x6501) );
CLKBUF_X2 inst_18864 ( .A(net_15643), .Z(net_18712) );
SDFF_X2 inst_768 ( .Q(net_8811), .D(net_8811), .SI(net_3976), .SE(net_3879), .CK(net_10525) );
SDFFR_X2 inst_2121 ( .SI(net_7185), .Q(net_7185), .D(net_6436), .SE(net_4362), .CK(net_13570), .RN(x6501) );
NAND2_X2 inst_4850 ( .ZN(net_1419), .A2(net_900), .A1(net_165) );
CLKBUF_X2 inst_12067 ( .A(net_11914), .Z(net_11915) );
INV_X16 inst_6639 ( .ZN(net_3934), .A(net_3336) );
CLKBUF_X2 inst_16450 ( .A(net_10180), .Z(net_16298) );
CLKBUF_X2 inst_11001 ( .A(net_10848), .Z(net_10849) );
CLKBUF_X2 inst_13225 ( .A(net_13072), .Z(net_13073) );
DFF_X1 inst_6774 ( .Q(net_7553), .D(net_4598), .CK(net_12761) );
NOR2_X2 inst_3494 ( .A1(net_8214), .ZN(net_2188), .A2(net_2187) );
CLKBUF_X2 inst_18960 ( .A(net_18807), .Z(net_18808) );
CLKBUF_X2 inst_17172 ( .A(net_17019), .Z(net_17020) );
SDFF_X2 inst_1867 ( .D(net_7268), .SI(net_6925), .Q(net_6925), .SE(net_6281), .CK(net_14340) );
CLKBUF_X2 inst_18997 ( .A(net_18844), .Z(net_18845) );
CLKBUF_X2 inst_17165 ( .A(net_13640), .Z(net_17013) );
CLKBUF_X2 inst_13627 ( .A(net_13474), .Z(net_13475) );
INV_X2 inst_6314 ( .ZN(net_3349), .A(net_3298) );
DFFR_X1 inst_7580 ( .D(net_6481), .Q(net_6463), .CK(net_15118), .RN(x6501) );
CLKBUF_X2 inst_18882 ( .A(net_18729), .Z(net_18730) );
DFFR_X2 inst_7046 ( .QN(net_8900), .D(net_4894), .CK(net_14496), .RN(x6501) );
CLKBUF_X2 inst_13782 ( .A(net_13629), .Z(net_13630) );
AOI22_X2 inst_7909 ( .B2(net_5609), .ZN(net_4516), .A2(net_4515), .A1(net_1655), .B1(net_382) );
INV_X4 inst_5670 ( .A(net_7488), .ZN(net_4699) );
CLKBUF_X2 inst_15222 ( .A(net_13964), .Z(net_15070) );
DFF_X1 inst_6791 ( .Q(net_8250), .D(net_4429), .CK(net_17605) );
CLKBUF_X2 inst_15862 ( .A(net_15709), .Z(net_15710) );
CLKBUF_X2 inst_13695 ( .A(net_13542), .Z(net_13543) );
CLKBUF_X2 inst_12575 ( .A(net_12422), .Z(net_12423) );
CLKBUF_X2 inst_14143 ( .A(net_13990), .Z(net_13991) );
NAND2_X1 inst_4912 ( .A1(net_6808), .A2(net_6805), .ZN(net_612) );
NOR2_X2 inst_3342 ( .A1(net_6337), .ZN(net_5939), .A2(net_5933) );
NAND2_X2 inst_4825 ( .ZN(net_1109), .A2(net_758), .A1(x4886) );
CLKBUF_X2 inst_9832 ( .A(net_9679), .Z(net_9680) );
CLKBUF_X2 inst_14666 ( .A(net_14513), .Z(net_14514) );
AOI22_X2 inst_8175 ( .B1(net_8863), .A1(net_8308), .B2(net_6252), .A2(net_4345), .ZN(net_3855) );
NAND3_X2 inst_3895 ( .ZN(net_5643), .A1(net_5572), .A3(net_5506), .A2(net_5414) );
XNOR2_X2 inst_303 ( .ZN(net_973), .A(net_972), .B(net_194) );
CLKBUF_X2 inst_13518 ( .A(net_13365), .Z(net_13366) );
CLKBUF_X2 inst_14324 ( .A(net_14171), .Z(net_14172) );
SDFF_X2 inst_1275 ( .Q(net_7809), .D(net_7809), .SE(net_2730), .SI(net_2655), .CK(net_15856) );
CLKBUF_X2 inst_18362 ( .A(net_18209), .Z(net_18210) );
XOR2_X2 inst_26 ( .Z(net_1357), .A(net_1356), .B(net_739) );
CLKBUF_X2 inst_15326 ( .A(net_15173), .Z(net_15174) );
CLKBUF_X2 inst_13052 ( .A(net_12899), .Z(net_12900) );
CLKBUF_X2 inst_10480 ( .A(net_9508), .Z(net_10328) );
AOI22_X2 inst_8104 ( .B1(net_8178), .A1(net_7736), .B2(net_6101), .A2(net_6095), .ZN(net_4044) );
CLKBUF_X2 inst_10198 ( .A(net_10045), .Z(net_10046) );
CLKBUF_X2 inst_17096 ( .A(net_16475), .Z(net_16944) );
CLKBUF_X2 inst_12731 ( .A(net_12578), .Z(net_12579) );
CLKBUF_X2 inst_14038 ( .A(net_13885), .Z(net_13886) );
CLKBUF_X2 inst_10001 ( .A(net_9848), .Z(net_9849) );
INV_X2 inst_6530 ( .A(net_6751), .ZN(net_522) );
DFFR_X1 inst_7490 ( .QN(net_6327), .D(net_3877), .CK(net_17645), .RN(x6501) );
CLKBUF_X2 inst_12895 ( .A(net_12742), .Z(net_12743) );
NAND2_X2 inst_4864 ( .A2(net_8269), .ZN(net_843), .A1(net_680) );
CLKBUF_X2 inst_15900 ( .A(net_15747), .Z(net_15748) );
CLKBUF_X2 inst_16211 ( .A(net_16058), .Z(net_16059) );
NAND4_X2 inst_3765 ( .ZN(net_4256), .A1(net_3797), .A2(net_3796), .A3(net_3795), .A4(net_3794) );
CLKBUF_X2 inst_15924 ( .A(net_15771), .Z(net_15772) );
CLKBUF_X2 inst_17056 ( .A(net_16903), .Z(net_16904) );
NAND2_X2 inst_4218 ( .A1(net_7013), .A2(net_5249), .ZN(net_5242) );
CLKBUF_X2 inst_15808 ( .A(net_15655), .Z(net_15656) );
CLKBUF_X2 inst_10062 ( .A(net_9200), .Z(net_9910) );
INV_X2 inst_6456 ( .A(net_7592), .ZN(net_3134) );
CLKBUF_X2 inst_16689 ( .A(net_16536), .Z(net_16537) );
CLKBUF_X2 inst_17511 ( .A(net_17358), .Z(net_17359) );
CLKBUF_X2 inst_16720 ( .A(net_16567), .Z(net_16568) );
DFFR_X2 inst_7064 ( .QN(net_7205), .D(net_4311), .CK(net_13598), .RN(x6501) );
CLKBUF_X2 inst_18020 ( .A(net_17867), .Z(net_17868) );
CLKBUF_X2 inst_11636 ( .A(net_11483), .Z(net_11484) );
CLKBUF_X2 inst_13702 ( .A(net_13549), .Z(net_13550) );
CLKBUF_X2 inst_11469 ( .A(net_10205), .Z(net_11317) );
INV_X8 inst_5053 ( .ZN(net_6253), .A(net_3376) );
CLKBUF_X2 inst_15137 ( .A(net_14984), .Z(net_14985) );
CLKBUF_X2 inst_18373 ( .A(net_11415), .Z(net_18221) );
CLKBUF_X2 inst_17484 ( .A(net_17331), .Z(net_17332) );
SDFF_X2 inst_1438 ( .SI(net_7282), .Q(net_7099), .D(net_7099), .SE(net_6278), .CK(net_14923) );
CLKBUF_X2 inst_10454 ( .A(net_10301), .Z(net_10302) );
INV_X2 inst_6373 ( .A(net_1739), .ZN(net_1595) );
CLKBUF_X2 inst_17795 ( .A(net_17642), .Z(net_17643) );
CLKBUF_X2 inst_18005 ( .A(net_17852), .Z(net_17853) );
CLKBUF_X2 inst_12681 ( .A(net_12528), .Z(net_12529) );
SDFF_X2 inst_880 ( .Q(net_8592), .D(net_8592), .SI(net_3948), .SE(net_3878), .CK(net_13463) );
CLKBUF_X2 inst_12241 ( .A(net_12088), .Z(net_12089) );
CLKBUF_X2 inst_11437 ( .A(net_11284), .Z(net_11285) );
CLKBUF_X2 inst_16596 ( .A(net_16443), .Z(net_16444) );
SDFFR_X1 inst_2681 ( .SI(net_7544), .SE(net_5043), .CK(net_9697), .RN(x6501), .Q(x4011), .D(x4011) );
NOR2_X2 inst_3445 ( .A1(net_6383), .A2(net_5902), .ZN(net_3114) );
AND2_X4 inst_9118 ( .ZN(net_1614), .A1(net_1467), .A2(net_1100) );
CLKBUF_X2 inst_12370 ( .A(net_12217), .Z(net_12218) );
CLKBUF_X2 inst_16023 ( .A(net_15870), .Z(net_15871) );
AND3_X4 inst_9044 ( .A2(net_2680), .ZN(net_2236), .A1(net_2077), .A3(net_1965) );
NAND3_X2 inst_3972 ( .ZN(net_2184), .A3(net_2183), .A1(net_1902), .A2(net_1316) );
HA_X1 inst_6670 ( .A(net_4457), .S(net_3223), .CO(net_3222), .B(net_3040) );
CLKBUF_X2 inst_11633 ( .A(net_11480), .Z(net_11481) );
CLKBUF_X2 inst_17186 ( .A(net_17033), .Z(net_17034) );
SDFF_X2 inst_1388 ( .SI(net_7293), .Q(net_7110), .D(net_7110), .SE(net_6278), .CK(net_18404) );
SDFFR_X1 inst_2699 ( .SI(net_7531), .SE(net_5043), .CK(net_11943), .RN(x6501), .Q(x4166), .D(x4166) );
NOR2_X2 inst_3517 ( .A2(net_3023), .ZN(net_1768), .A1(net_1449) );
CLKBUF_X2 inst_9291 ( .A(net_9138), .Z(net_9139) );
CLKBUF_X2 inst_14927 ( .A(net_13198), .Z(net_14775) );
AOI22_X2 inst_8506 ( .B1(net_6654), .A1(net_6621), .A2(net_6213), .B2(net_6138), .ZN(net_3434) );
NOR2_X2 inst_3396 ( .ZN(net_4537), .A1(net_4371), .A2(net_4370) );
SDFF_X2 inst_1372 ( .Q(net_8182), .D(net_8182), .SI(net_2705), .SE(net_2561), .CK(net_18552) );
DFFR_X2 inst_7332 ( .D(net_7627), .Q(net_7618), .CK(net_17986), .RN(x6501) );
CLKBUF_X2 inst_12109 ( .A(net_11956), .Z(net_11957) );
CLKBUF_X2 inst_10631 ( .A(net_10478), .Z(net_10479) );
CLKBUF_X2 inst_9759 ( .A(net_9606), .Z(net_9607) );
INV_X4 inst_6081 ( .A(net_7164), .ZN(net_835) );
SDFFR_X1 inst_2761 ( .QN(net_7593), .SE(net_3144), .SI(net_2836), .D(net_1497), .CK(net_13453), .RN(x6501) );
SDFF_X2 inst_989 ( .D(net_7327), .SI(net_6635), .Q(net_6635), .SE(net_3123), .CK(net_11333) );
CLKBUF_X2 inst_15087 ( .A(net_14934), .Z(net_14935) );
SDFFR_X2 inst_2283 ( .SI(net_7396), .SE(net_2789), .Q(net_255), .D(net_255), .CK(net_18329), .RN(x6501) );
SDFF_X2 inst_858 ( .Q(net_8556), .D(net_8556), .SI(net_3961), .SE(net_3878), .CK(net_13165) );
CLKBUF_X2 inst_19080 ( .A(net_18722), .Z(net_18928) );
AND2_X4 inst_9111 ( .ZN(net_2037), .A2(net_1849), .A1(net_521) );
CLKBUF_X2 inst_13779 ( .A(net_11793), .Z(net_13627) );
CLKBUF_X2 inst_12060 ( .A(net_11907), .Z(net_11908) );
OAI22_X2 inst_2936 ( .ZN(net_2045), .A1(net_2043), .B1(net_1858), .A2(net_1790), .B2(net_1136) );
SDFFR_X2 inst_2468 ( .D(net_4714), .SE(net_2757), .SI(net_409), .Q(net_409), .CK(net_16651), .RN(x6501) );
XOR2_X2 inst_54 ( .A(net_3533), .Z(net_993), .B(net_551) );
CLKBUF_X2 inst_12610 ( .A(net_12457), .Z(net_12458) );
CLKBUF_X2 inst_10556 ( .A(net_10340), .Z(net_10404) );
SDFF_X2 inst_1482 ( .SI(net_7271), .Q(net_7048), .D(net_7048), .SE(net_6280), .CK(net_16831) );
SDFF_X2 inst_1420 ( .SI(net_7266), .Q(net_7043), .D(net_7043), .SE(net_6280), .CK(net_17091) );
CLKBUF_X2 inst_18678 ( .A(net_18525), .Z(net_18526) );
CLKBUF_X2 inst_12177 ( .A(net_12024), .Z(net_12025) );
CLKBUF_X2 inst_12988 ( .A(net_12835), .Z(net_12836) );
INV_X4 inst_5337 ( .ZN(net_1593), .A(net_1458) );
NAND2_X2 inst_4062 ( .ZN(net_5879), .A2(net_5769), .A1(net_3280) );
INV_X4 inst_5730 ( .A(net_7238), .ZN(net_1956) );
CLKBUF_X2 inst_16819 ( .A(net_16666), .Z(net_16667) );
CLKBUF_X2 inst_15775 ( .A(net_15622), .Z(net_15623) );
CLKBUF_X2 inst_15685 ( .A(net_15532), .Z(net_15533) );
NAND2_X2 inst_4108 ( .ZN(net_5423), .A2(net_5238), .A1(net_5147) );
NAND2_X2 inst_4626 ( .A2(net_2835), .ZN(net_2834), .A1(net_1739) );
AOI221_X2 inst_8780 ( .B1(net_7187), .C2(net_6187), .B2(net_5655), .ZN(net_5258), .A(net_4934), .C1(net_188) );
CLKBUF_X2 inst_9491 ( .A(net_9338), .Z(net_9339) );
CLKBUF_X2 inst_11595 ( .A(net_11442), .Z(net_11443) );
CLKBUF_X2 inst_15496 ( .A(net_15343), .Z(net_15344) );
CLKBUF_X2 inst_15272 ( .A(net_15119), .Z(net_15120) );
SDFF_X2 inst_497 ( .SI(net_8595), .Q(net_8595), .SE(net_3984), .D(net_3980), .CK(net_10738) );
CLKBUF_X2 inst_13826 ( .A(net_13673), .Z(net_13674) );
DFFR_X1 inst_7517 ( .Q(net_7216), .D(net_1602), .CK(net_18968), .RN(x6501) );
CLKBUF_X2 inst_18320 ( .A(net_18167), .Z(net_18168) );
CLKBUF_X2 inst_15919 ( .A(net_14818), .Z(net_15767) );
SDFFR_X2 inst_2195 ( .QN(net_7224), .SI(net_2931), .D(net_2665), .SE(net_1379), .CK(net_15147), .RN(x6501) );
AOI221_X2 inst_8787 ( .B2(net_6450), .B1(net_5654), .C2(net_5595), .ZN(net_5023), .A(net_5022), .C1(net_332) );
SDFF_X2 inst_1335 ( .SI(net_7681), .Q(net_7681), .SE(net_2714), .D(net_2706), .CK(net_18078) );
CLKBUF_X2 inst_15197 ( .A(net_12040), .Z(net_15045) );
CLKBUF_X2 inst_9924 ( .A(net_9771), .Z(net_9772) );
NAND4_X2 inst_3845 ( .ZN(net_1698), .A2(net_1426), .A1(net_1412), .A3(net_1410), .A4(net_1400) );
DFFR_X2 inst_7173 ( .QN(net_7349), .D(net_2799), .CK(net_9566), .RN(x6501) );
CLKBUF_X2 inst_10124 ( .A(net_9162), .Z(net_9972) );
INV_X4 inst_5168 ( .ZN(net_3027), .A(net_3026) );
OAI21_X2 inst_3128 ( .ZN(net_2211), .B1(net_2159), .B2(net_2157), .A(net_1098) );
CLKBUF_X2 inst_10715 ( .A(net_10562), .Z(net_10563) );
CLKBUF_X2 inst_17749 ( .A(net_12755), .Z(net_17597) );
CLKBUF_X2 inst_14653 ( .A(net_14500), .Z(net_14501) );
SDFFR_X2 inst_2517 ( .D(net_7392), .SE(net_2378), .SI(net_225), .Q(net_225), .CK(net_17753), .RN(x6501) );
NAND2_X2 inst_4183 ( .ZN(net_5320), .A1(net_5074), .A2(net_5073) );
CLKBUF_X2 inst_10806 ( .A(net_10653), .Z(net_10654) );
SDFF_X2 inst_714 ( .SI(net_8659), .Q(net_8659), .D(net_3952), .SE(net_3885), .CK(net_12876) );
CLKBUF_X2 inst_15735 ( .A(net_15041), .Z(net_15583) );
CLKBUF_X2 inst_15518 ( .A(net_15365), .Z(net_15366) );
OAI21_X2 inst_3005 ( .ZN(net_5761), .A(net_5756), .B2(net_5755), .B1(net_660) );
OR2_X2 inst_2895 ( .ZN(net_1289), .A2(net_1063), .A1(net_638) );
AOI211_X2 inst_9005 ( .C2(net_5657), .ZN(net_5584), .B(net_5285), .A(net_4825), .C1(net_509) );
CLKBUF_X2 inst_16199 ( .A(net_16046), .Z(net_16047) );
SDFF_X2 inst_1061 ( .D(net_7333), .SI(net_6641), .Q(net_6641), .SE(net_3123), .CK(net_11681) );
CLKBUF_X2 inst_11201 ( .A(net_11048), .Z(net_11049) );
SDFFR_X2 inst_2326 ( .SE(net_2260), .Q(net_371), .D(net_371), .CK(net_11393), .RN(x6501), .SI(x1639) );
INV_X1 inst_6657 ( .A(net_6183), .ZN(net_6180) );
CLKBUF_X2 inst_18183 ( .A(net_14030), .Z(net_18031) );
XOR2_X1 inst_72 ( .Z(net_3391), .B(net_3390), .A(net_3228) );
DFFR_X2 inst_6967 ( .QN(net_6343), .D(net_5939), .CK(net_17484), .RN(x6501) );
CLKBUF_X2 inst_11703 ( .A(net_11550), .Z(net_11551) );
CLKBUF_X2 inst_17920 ( .A(net_17767), .Z(net_17768) );
SDFF_X2 inst_1634 ( .Q(net_8179), .D(net_8179), .SI(net_2703), .SE(net_2538), .CK(net_14006) );
CLKBUF_X2 inst_15961 ( .A(net_12464), .Z(net_15809) );
AOI21_X2 inst_8998 ( .ZN(net_1305), .B2(net_1304), .B1(x13208), .A(x13193) );
AOI22_X2 inst_7980 ( .B1(net_8027), .A1(net_7993), .B2(net_6102), .A2(net_6097), .ZN(net_6038) );
CLKBUF_X2 inst_10619 ( .A(net_10260), .Z(net_10467) );
DFF_X1 inst_6729 ( .Q(net_6756), .D(net_5640), .CK(net_10444) );
INV_X16 inst_6650 ( .ZN(net_6190), .A(net_4415) );
CLKBUF_X2 inst_19114 ( .A(net_18951), .Z(net_18962) );
CLKBUF_X2 inst_15609 ( .A(net_15456), .Z(net_15457) );
CLKBUF_X2 inst_9485 ( .A(net_9332), .Z(net_9333) );
CLKBUF_X2 inst_12415 ( .A(net_12262), .Z(net_12263) );
CLKBUF_X2 inst_12357 ( .A(net_10483), .Z(net_12205) );
NAND2_X2 inst_4638 ( .ZN(net_2442), .A2(net_2440), .A1(net_2344) );
CLKBUF_X2 inst_11487 ( .A(net_11334), .Z(net_11335) );
CLKBUF_X2 inst_13426 ( .A(net_10286), .Z(net_13274) );
SDFF_X2 inst_1582 ( .Q(net_8035), .D(net_8035), .SI(net_2711), .SE(net_2545), .CK(net_17069) );
CLKBUF_X2 inst_16122 ( .A(net_11006), .Z(net_15970) );
CLKBUF_X2 inst_13202 ( .A(net_12422), .Z(net_13050) );
CLKBUF_X2 inst_17585 ( .A(net_17432), .Z(net_17433) );
INV_X2 inst_6334 ( .ZN(net_2900), .A(net_2899) );
CLKBUF_X2 inst_13905 ( .A(net_13395), .Z(net_13753) );
INV_X4 inst_5846 ( .A(net_6388), .ZN(net_1188) );
CLKBUF_X2 inst_18858 ( .A(net_18705), .Z(net_18706) );
SDFF_X2 inst_1840 ( .D(net_7287), .SI(net_6904), .Q(net_6904), .SE(net_6284), .CK(net_14891) );
INV_X2 inst_6345 ( .ZN(net_2444), .A(net_2443) );
XNOR2_X2 inst_133 ( .B(net_6404), .ZN(net_2813), .A(net_2465) );
CLKBUF_X2 inst_17805 ( .A(net_17652), .Z(net_17653) );
CLKBUF_X2 inst_14734 ( .A(net_10129), .Z(net_14582) );
CLKBUF_X2 inst_13847 ( .A(net_10109), .Z(net_13695) );
CLKBUF_X2 inst_16587 ( .A(net_16434), .Z(net_16435) );
CLKBUF_X2 inst_18955 ( .A(net_16771), .Z(net_18803) );
CLKBUF_X2 inst_9988 ( .A(net_9588), .Z(net_9836) );
CLKBUF_X2 inst_18552 ( .A(net_18399), .Z(net_18400) );
CLKBUF_X2 inst_14688 ( .A(net_14535), .Z(net_14536) );
SDFF_X2 inst_1721 ( .Q(net_8117), .D(net_8117), .SI(net_2659), .SE(net_2541), .CK(net_15494) );
CLKBUF_X2 inst_9744 ( .A(net_9591), .Z(net_9592) );
CLKBUF_X2 inst_10884 ( .A(net_10731), .Z(net_10732) );
CLKBUF_X2 inst_18930 ( .A(net_17196), .Z(net_18778) );
CLKBUF_X2 inst_12854 ( .A(net_12701), .Z(net_12702) );
XNOR2_X2 inst_126 ( .ZN(net_2867), .B(net_2810), .A(net_2809) );
CLKBUF_X2 inst_18413 ( .A(net_18260), .Z(net_18261) );
NAND3_X2 inst_3887 ( .ZN(net_5651), .A1(net_5580), .A3(net_5514), .A2(net_5448) );
CLKBUF_X2 inst_14163 ( .A(net_12553), .Z(net_14011) );
SDFF_X2 inst_1631 ( .Q(net_8148), .D(net_8148), .SI(net_2705), .SE(net_2538), .CK(net_18549) );
CLKBUF_X2 inst_12651 ( .A(net_12220), .Z(net_12499) );
DFFR_X1 inst_7510 ( .D(net_1686), .Q(net_390), .CK(net_13539), .RN(x6501) );
CLKBUF_X2 inst_13106 ( .A(net_12953), .Z(net_12954) );
SDFF_X2 inst_1086 ( .D(net_7340), .SI(net_6516), .Q(net_6516), .SE(net_3071), .CK(net_11883) );
CLKBUF_X2 inst_14360 ( .A(net_14207), .Z(net_14208) );
SDFFR_X1 inst_2643 ( .D(net_6766), .SE(net_4506), .CK(net_9334), .RN(x6501), .SI(x1885), .Q(x1885) );
CLKBUF_X2 inst_12088 ( .A(net_11935), .Z(net_11936) );
CLKBUF_X2 inst_18354 ( .A(net_18201), .Z(net_18202) );
CLKBUF_X2 inst_13950 ( .A(net_10382), .Z(net_13798) );
CLKBUF_X2 inst_12615 ( .A(net_12462), .Z(net_12463) );
CLKBUF_X2 inst_12713 ( .A(net_12560), .Z(net_12561) );
SDFF_X2 inst_1688 ( .Q(net_8158), .D(net_8158), .SI(net_2574), .SE(net_2538), .CK(net_16033) );
CLKBUF_X2 inst_15621 ( .A(net_15468), .Z(net_15469) );
CLKBUF_X2 inst_13651 ( .A(net_13498), .Z(net_13499) );
CLKBUF_X2 inst_13732 ( .A(net_9576), .Z(net_13580) );
CLKBUF_X2 inst_17481 ( .A(net_10439), .Z(net_17329) );
CLKBUF_X2 inst_12146 ( .A(net_10935), .Z(net_11994) );
CLKBUF_X2 inst_14836 ( .A(net_14683), .Z(net_14684) );
CLKBUF_X2 inst_17580 ( .A(net_17427), .Z(net_17428) );
CLKBUF_X2 inst_13084 ( .A(net_12931), .Z(net_12932) );
SDFF_X2 inst_914 ( .SI(net_8706), .Q(net_8706), .SE(net_6195), .D(net_3980), .CK(net_10683) );
INV_X2 inst_6364 ( .A(net_2159), .ZN(net_1966) );
INV_X4 inst_5170 ( .ZN(net_3146), .A(net_3144) );
INV_X4 inst_5182 ( .ZN(net_2940), .A(net_2844) );
CLKBUF_X2 inst_12198 ( .A(net_12045), .Z(net_12046) );
CLKBUF_X2 inst_14962 ( .A(net_14809), .Z(net_14810) );
CLKBUF_X2 inst_11588 ( .A(net_10548), .Z(net_11436) );
SDFF_X2 inst_384 ( .SI(net_8384), .Q(net_8384), .SE(net_3969), .D(net_3966), .CK(net_10040) );
SDFF_X2 inst_1252 ( .SI(net_7698), .Q(net_7698), .D(net_2715), .SE(net_2714), .CK(net_16874) );
CLKBUF_X2 inst_12773 ( .A(net_12620), .Z(net_12621) );
NAND4_X2 inst_3800 ( .ZN(net_3626), .A1(net_3487), .A2(net_3486), .A3(net_3485), .A4(net_3484) );
CLKBUF_X2 inst_17568 ( .A(net_14403), .Z(net_17416) );
CLKBUF_X2 inst_17458 ( .A(net_17204), .Z(net_17306) );
INV_X4 inst_6086 ( .A(net_6293), .ZN(net_2670) );
CLKBUF_X2 inst_12989 ( .A(net_9337), .Z(net_12837) );
CLKBUF_X2 inst_10271 ( .A(net_10063), .Z(net_10119) );
SDFFR_X2 inst_2209 ( .Q(net_8942), .D(net_2472), .SI(net_1991), .SE(net_1474), .CK(net_16258), .RN(x6501) );
SDFFR_X1 inst_2722 ( .SI(net_9032), .Q(net_9032), .D(net_7461), .SE(net_3208), .CK(net_10669), .RN(x6501) );
CLKBUF_X2 inst_13034 ( .A(net_12881), .Z(net_12882) );
CLKBUF_X2 inst_17738 ( .A(net_17585), .Z(net_17586) );
CLKBUF_X2 inst_19093 ( .A(net_18940), .Z(net_18941) );
CLKBUF_X2 inst_16817 ( .A(net_16664), .Z(net_16665) );
SDFF_X2 inst_1238 ( .Q(net_7957), .D(net_7957), .SE(net_2755), .SI(net_2576), .CK(net_16009) );
DFFR_X2 inst_7361 ( .Q(net_7341), .CK(net_11706), .D(x12902), .RN(x6501) );
SDFFR_X2 inst_2171 ( .QN(net_7569), .D(net_3937), .SE(net_3144), .SI(net_3130), .CK(net_13077), .RN(x6501) );
CLKBUF_X2 inst_15385 ( .A(net_15232), .Z(net_15233) );
AND4_X4 inst_9031 ( .A3(net_8960), .ZN(net_1670), .A2(net_1334), .A4(net_1169), .A1(net_910) );
AOI22_X2 inst_7941 ( .B1(net_8123), .A1(net_7885), .A2(net_6098), .B2(net_4190), .ZN(net_4184) );
AOI22_X2 inst_8527 ( .B1(net_6590), .A1(net_6557), .A2(net_6257), .B2(net_6110), .ZN(net_3413) );
NOR2_X2 inst_3402 ( .A2(net_6424), .ZN(net_4401), .A1(net_2849) );
CLKBUF_X2 inst_18616 ( .A(net_18463), .Z(net_18464) );
CLKBUF_X2 inst_14318 ( .A(net_14165), .Z(net_14166) );
SDFF_X2 inst_1011 ( .SI(net_7324), .Q(net_6665), .D(net_6665), .SE(net_3126), .CK(net_9870) );
SDFF_X2 inst_404 ( .SI(net_8317), .Q(net_8317), .SE(net_3978), .D(net_3957), .CK(net_13295) );
INV_X4 inst_5838 ( .A(net_8892), .ZN(net_3000) );
NOR2_X2 inst_3615 ( .ZN(net_1062), .A2(x12810), .A1(x12780) );
CLKBUF_X2 inst_9628 ( .A(net_9475), .Z(net_9476) );
OAI211_X2 inst_3216 ( .ZN(net_3023), .C2(net_1802), .C1(net_1723), .B(net_1631), .A(net_1513) );
AOI221_X2 inst_8748 ( .B2(net_5657), .ZN(net_5610), .C2(net_5609), .A(net_5517), .B1(net_2694), .C1(net_364) );
CLKBUF_X2 inst_15093 ( .A(net_14940), .Z(net_14941) );
CLKBUF_X2 inst_18228 ( .A(net_18075), .Z(net_18076) );
CLKBUF_X2 inst_15489 ( .A(net_15336), .Z(net_15337) );
NOR2_X2 inst_3540 ( .ZN(net_2269), .A1(net_1452), .A2(net_1130) );
CLKBUF_X2 inst_15277 ( .A(net_15124), .Z(net_15125) );
CLKBUF_X2 inst_17723 ( .A(net_15577), .Z(net_17571) );
CLKBUF_X2 inst_14005 ( .A(net_13852), .Z(net_13853) );
CLKBUF_X2 inst_10904 ( .A(net_9295), .Z(net_10752) );
CLKBUF_X2 inst_18541 ( .A(net_12076), .Z(net_18389) );
SDFFR_X2 inst_2413 ( .SE(net_2748), .D(net_630), .SI(net_455), .Q(net_455), .CK(net_13948), .RN(x6501) );
SDFF_X2 inst_1574 ( .Q(net_8024), .D(net_8024), .SI(net_2589), .SE(net_2545), .CK(net_15268) );
CLKBUF_X2 inst_18755 ( .A(net_18602), .Z(net_18603) );
CLKBUF_X2 inst_16549 ( .A(net_16396), .Z(net_16397) );
DFFR_X1 inst_7528 ( .Q(net_7660), .D(net_7656), .CK(net_12718), .RN(x6501) );
CLKBUF_X2 inst_14518 ( .A(net_14365), .Z(net_14366) );
XNOR2_X2 inst_228 ( .A(net_3082), .ZN(net_1358), .B(net_1356) );
CLKBUF_X2 inst_14034 ( .A(net_13881), .Z(net_13882) );
DFFS_X2 inst_6872 ( .Q(net_8895), .D(net_3971), .CK(net_11203), .SN(x6501) );
CLKBUF_X2 inst_12008 ( .A(net_11713), .Z(net_11856) );
CLKBUF_X2 inst_19019 ( .A(net_13092), .Z(net_18867) );
CLKBUF_X2 inst_12279 ( .A(net_9326), .Z(net_12127) );
AOI221_X2 inst_8759 ( .C2(net_6130), .B2(net_5535), .ZN(net_5473), .A(net_4953), .C1(net_1381), .B1(net_465) );
XNOR2_X2 inst_244 ( .B(net_6821), .ZN(net_1217), .A(net_1216) );
CLKBUF_X2 inst_18801 ( .A(net_18648), .Z(net_18649) );
CLKBUF_X2 inst_17881 ( .A(net_13157), .Z(net_17729) );
CLKBUF_X2 inst_13514 ( .A(net_10444), .Z(net_13362) );
INV_X4 inst_5262 ( .A(net_1771), .ZN(net_1770) );
CLKBUF_X2 inst_11472 ( .A(net_11319), .Z(net_11320) );
CLKBUF_X2 inst_13464 ( .A(net_13311), .Z(net_13312) );
CLKBUF_X2 inst_12136 ( .A(net_11983), .Z(net_11984) );
CLKBUF_X2 inst_11794 ( .A(net_11641), .Z(net_11642) );
INV_X4 inst_5537 ( .ZN(net_1175), .A(net_742) );
CLKBUF_X2 inst_18887 ( .A(net_15614), .Z(net_18735) );
CLKBUF_X2 inst_11339 ( .A(net_10468), .Z(net_11187) );
OAI21_X2 inst_3079 ( .ZN(net_3536), .A(net_3535), .B1(net_3311), .B2(net_3300) );
CLKBUF_X2 inst_16951 ( .A(net_16798), .Z(net_16799) );
CLKBUF_X2 inst_10143 ( .A(net_9066), .Z(net_9991) );
CLKBUF_X2 inst_12529 ( .A(net_12376), .Z(net_12377) );
INV_X4 inst_5487 ( .A(net_1994), .ZN(net_729) );
CLKBUF_X2 inst_11789 ( .A(net_11636), .Z(net_11637) );
CLKBUF_X2 inst_10303 ( .A(net_10150), .Z(net_10151) );
CLKBUF_X2 inst_18949 ( .A(net_18796), .Z(net_18797) );
NOR2_X2 inst_3606 ( .A2(net_1757), .A1(net_1450), .ZN(net_1334) );
XOR2_X1 inst_93 ( .Z(net_1416), .B(net_1415), .A(net_621) );
CLKBUF_X2 inst_17192 ( .A(net_17039), .Z(net_17040) );
NAND2_X2 inst_4832 ( .A2(net_5957), .ZN(net_1812), .A1(net_601) );
DFFR_X2 inst_7026 ( .QN(net_6289), .D(net_5685), .CK(net_13867), .RN(x6501) );
CLKBUF_X2 inst_14631 ( .A(net_14478), .Z(net_14479) );
CLKBUF_X2 inst_17632 ( .A(net_9750), .Z(net_17480) );
CLKBUF_X2 inst_12105 ( .A(net_11952), .Z(net_11953) );
AOI22_X2 inst_7784 ( .A1(net_5268), .ZN(net_4866), .A2(net_4631), .B2(net_4388), .B1(net_2628) );
NAND2_X2 inst_4595 ( .A2(net_6407), .ZN(net_2908), .A1(net_2530) );
SDFF_X2 inst_1675 ( .SI(net_7744), .Q(net_7744), .D(net_2708), .SE(net_2560), .CK(net_15501) );
CLKBUF_X2 inst_11086 ( .A(net_9539), .Z(net_10934) );
NOR2_X2 inst_3433 ( .A2(net_3093), .ZN(net_3076), .A1(net_1672) );
CLKBUF_X2 inst_11274 ( .A(net_9457), .Z(net_11122) );
INV_X4 inst_5149 ( .ZN(net_3243), .A(net_3211) );
AOI21_X2 inst_8958 ( .ZN(net_4867), .A(net_4683), .B2(net_4564), .B1(net_232) );
CLKBUF_X2 inst_13713 ( .A(net_9858), .Z(net_13561) );
NAND2_X2 inst_4237 ( .A1(net_6901), .A2(net_5247), .ZN(net_5223) );
CLKBUF_X2 inst_10709 ( .A(net_10051), .Z(net_10557) );
XNOR2_X2 inst_148 ( .ZN(net_2117), .A(net_1839), .B(net_1827) );
SDFF_X2 inst_554 ( .Q(net_8701), .D(net_8701), .SI(net_3939), .SE(net_3935), .CK(net_11013) );
CLKBUF_X2 inst_13675 ( .A(net_9459), .Z(net_13523) );
CLKBUF_X2 inst_13621 ( .A(net_12399), .Z(net_13469) );
SDFF_X2 inst_1187 ( .D(net_7342), .SI(net_6584), .Q(net_6584), .SE(net_3070), .CK(net_9439) );
INV_X4 inst_6000 ( .A(net_8959), .ZN(net_1846) );
INV_X4 inst_5499 ( .ZN(net_704), .A(net_703) );
CLKBUF_X2 inst_19147 ( .A(net_18994), .Z(net_18995) );
CLKBUF_X2 inst_17963 ( .A(net_17810), .Z(net_17811) );
CLKBUF_X2 inst_10740 ( .A(net_10587), .Z(net_10588) );
AOI21_X2 inst_8951 ( .A(net_5783), .ZN(net_5666), .B1(net_5470), .B2(net_5264) );
SDFF_X2 inst_1917 ( .D(net_7268), .SI(net_6845), .Q(net_6845), .SE(net_6282), .CK(net_14329) );
CLKBUF_X2 inst_14764 ( .A(net_14611), .Z(net_14612) );
CLKBUF_X2 inst_19060 ( .A(net_10114), .Z(net_18908) );
CLKBUF_X2 inst_15302 ( .A(net_10087), .Z(net_15150) );
CLKBUF_X2 inst_15753 ( .A(net_15600), .Z(net_15601) );
CLKBUF_X2 inst_12695 ( .A(net_12542), .Z(net_12543) );
MUX2_X2 inst_4955 ( .A(net_7380), .S(net_2376), .Z(net_2368), .B(net_886) );
CLKBUF_X2 inst_11553 ( .A(net_11400), .Z(net_11401) );
CLKBUF_X2 inst_12386 ( .A(net_9110), .Z(net_12234) );
CLKBUF_X2 inst_16292 ( .A(net_16139), .Z(net_16140) );
CLKBUF_X2 inst_17909 ( .A(net_10288), .Z(net_17757) );
SDFFS_X2 inst_2087 ( .SI(net_6344), .SE(net_1136), .CK(net_16526), .SN(x6501), .Q(x971), .D(x971) );
CLKBUF_X2 inst_16215 ( .A(net_16062), .Z(net_16063) );
CLKBUF_X2 inst_13891 ( .A(net_13738), .Z(net_13739) );
CLKBUF_X2 inst_15671 ( .A(net_15518), .Z(net_15519) );
CLKBUF_X2 inst_19058 ( .A(net_18905), .Z(net_18906) );
CLKBUF_X2 inst_9881 ( .A(net_9258), .Z(net_9729) );
AOI22_X2 inst_8571 ( .B1(net_8941), .A1(net_8254), .B2(net_6164), .A2(net_6161), .ZN(net_2003) );
CLKBUF_X2 inst_16858 ( .A(net_16705), .Z(net_16706) );
INV_X2 inst_6501 ( .A(net_5952), .ZN(net_897) );
SDFF_X2 inst_819 ( .SI(net_8511), .Q(net_8511), .D(net_3952), .SE(net_3884), .CK(net_10327) );
NAND2_X2 inst_4464 ( .ZN(net_4784), .A2(net_4783), .A1(x1195) );
NOR3_X2 inst_3320 ( .A3(net_7305), .ZN(net_1264), .A1(net_1237), .A2(net_821) );
SDFF_X2 inst_1468 ( .SI(net_7293), .Q(net_7150), .D(net_7150), .SE(net_6279), .CK(net_18398) );
CLKBUF_X2 inst_9663 ( .A(net_9184), .Z(net_9511) );
CLKBUF_X2 inst_18068 ( .A(net_17915), .Z(net_17916) );
NAND4_X2 inst_3776 ( .ZN(net_4245), .A1(net_3730), .A2(net_3729), .A3(net_3728), .A4(net_3727) );
CLKBUF_X2 inst_18244 ( .A(net_18091), .Z(net_18092) );
CLKBUF_X2 inst_14046 ( .A(net_13893), .Z(net_13894) );
CLKBUF_X2 inst_16992 ( .A(net_16839), .Z(net_16840) );
AOI221_X2 inst_8857 ( .B1(net_8562), .C1(net_8451), .C2(net_6263), .B2(net_6262), .ZN(net_6233), .A(net_4234) );
INV_X4 inst_5859 ( .A(net_6396), .ZN(net_2494) );
CLKBUF_X2 inst_17641 ( .A(net_17488), .Z(net_17489) );
SDFFR_X2 inst_2617 ( .Q(net_7373), .D(net_7373), .SE(net_1136), .CK(net_18633), .RN(x6501), .SI(x4796) );
NAND3_X2 inst_3942 ( .A3(net_6328), .ZN(net_5679), .A2(net_4402), .A1(net_1702) );
CLKBUF_X2 inst_9459 ( .A(net_9306), .Z(net_9307) );
OAI21_X2 inst_3068 ( .B2(net_6425), .B1(net_4362), .ZN(net_4313), .A(net_2958) );
INV_X4 inst_5850 ( .A(net_7390), .ZN(net_1776) );
CLKBUF_X2 inst_18716 ( .A(net_16745), .Z(net_18564) );
SDFFR_X2 inst_2277 ( .SI(net_7390), .SE(net_2789), .Q(net_249), .D(net_249), .CK(net_14964), .RN(x6501) );
CLKBUF_X2 inst_9518 ( .A(net_9365), .Z(net_9366) );
CLKBUF_X2 inst_18335 ( .A(net_14349), .Z(net_18183) );
AOI22_X2 inst_8245 ( .B1(net_8576), .A1(net_8465), .A2(net_6263), .B2(net_6262), .ZN(net_3792) );
OAI221_X2 inst_2962 ( .C1(net_6752), .B1(net_6460), .ZN(net_3338), .B2(net_3174), .C2(net_3122), .A(net_3121) );
CLKBUF_X2 inst_16455 ( .A(net_16302), .Z(net_16303) );
CLKBUF_X2 inst_18940 ( .A(net_11163), .Z(net_18788) );
CLKBUF_X2 inst_13973 ( .A(net_13820), .Z(net_13821) );
CLKBUF_X2 inst_10605 ( .A(net_10452), .Z(net_10453) );
CLKBUF_X2 inst_9973 ( .A(net_9820), .Z(net_9821) );
XNOR2_X2 inst_208 ( .B(net_4699), .ZN(net_1485), .A(net_1484) );
CLKBUF_X2 inst_13756 ( .A(net_13603), .Z(net_13604) );
CLKBUF_X2 inst_16477 ( .A(net_16324), .Z(net_16325) );
CLKBUF_X2 inst_14272 ( .A(net_14119), .Z(net_14120) );
CLKBUF_X2 inst_15247 ( .A(net_15094), .Z(net_15095) );
NAND2_X2 inst_4202 ( .ZN(net_5294), .A1(net_5175), .A2(net_4980) );
NAND4_X2 inst_3774 ( .A3(net_6069), .A1(net_6068), .ZN(net_4247), .A2(net_3742), .A4(net_3741) );
DFFR_X2 inst_7101 ( .QN(net_7350), .D(net_3256), .CK(net_9570), .RN(x6501) );
INV_X4 inst_5282 ( .ZN(net_1630), .A(net_1531) );
CLKBUF_X2 inst_12751 ( .A(net_9465), .Z(net_12599) );
CLKBUF_X2 inst_11935 ( .A(net_11782), .Z(net_11783) );
CLKBUF_X2 inst_10294 ( .A(net_10141), .Z(net_10142) );
SDFF_X2 inst_636 ( .SI(net_8550), .Q(net_8550), .SE(net_3979), .D(net_3951), .CK(net_10599) );
CLKBUF_X2 inst_15823 ( .A(net_14476), .Z(net_15671) );
CLKBUF_X2 inst_18868 ( .A(net_18715), .Z(net_18716) );
CLKBUF_X2 inst_12499 ( .A(net_12346), .Z(net_12347) );
CLKBUF_X2 inst_11777 ( .A(net_11624), .Z(net_11625) );
CLKBUF_X2 inst_17208 ( .A(net_14168), .Z(net_17056) );
SDFF_X2 inst_1907 ( .D(net_7271), .SI(net_7008), .Q(net_7008), .SE(net_6277), .CK(net_16797) );
DFFR_X2 inst_7015 ( .QN(net_6296), .D(net_5741), .CK(net_16737), .RN(x6501) );
AOI22_X2 inst_8384 ( .B1(net_8746), .A1(net_8376), .A2(net_3867), .B2(net_3866), .ZN(net_3664) );
CLKBUF_X2 inst_16672 ( .A(net_16519), .Z(net_16520) );
CLKBUF_X2 inst_17859 ( .A(net_17706), .Z(net_17707) );
CLKBUF_X2 inst_10313 ( .A(net_10160), .Z(net_10161) );
CLKBUF_X2 inst_17169 ( .A(net_17016), .Z(net_17017) );
NAND4_X2 inst_3836 ( .A3(net_7524), .A1(net_4926), .ZN(net_2098), .A4(net_2097), .A2(net_1815) );
DFFR_X2 inst_6999 ( .QN(net_5967), .D(net_5882), .CK(net_9279), .RN(x6501) );
CLKBUF_X2 inst_13461 ( .A(net_13308), .Z(net_13309) );
AOI22_X2 inst_8472 ( .B1(net_6541), .A1(net_6508), .A2(net_6137), .B2(net_6104), .ZN(net_3468) );
SDFFR_X2 inst_2192 ( .SE(net_2588), .D(net_2587), .SI(net_385), .Q(net_385), .CK(net_10784), .RN(x6501) );
INV_X4 inst_5980 ( .A(net_5962), .ZN(x2948) );
AOI22_X2 inst_7806 ( .A2(net_8226), .A1(net_5268), .ZN(net_4768), .B1(net_4736), .B2(net_4388) );
CLKBUF_X2 inst_14675 ( .A(net_14522), .Z(net_14523) );
NAND2_X2 inst_4216 ( .A1(net_7012), .A2(net_5249), .ZN(net_5244) );
XOR2_X1 inst_106 ( .A(net_6817), .Z(net_992), .B(net_527) );
SDFFR_X2 inst_2583 ( .QN(net_7251), .D(net_2796), .SI(net_1954), .SE(net_1379), .CK(net_15350), .RN(x6501) );
CLKBUF_X2 inst_10753 ( .A(net_10600), .Z(net_10601) );
NAND3_X2 inst_3997 ( .A2(net_2981), .A1(net_1618), .ZN(net_1605), .A3(net_1499) );
CLKBUF_X2 inst_11344 ( .A(net_11191), .Z(net_11192) );
CLKBUF_X2 inst_16685 ( .A(net_16532), .Z(net_16533) );
INV_X4 inst_5241 ( .A(net_7299), .ZN(net_2544) );
CLKBUF_X2 inst_9903 ( .A(net_9245), .Z(net_9751) );
NAND2_X2 inst_4383 ( .A1(net_7158), .A2(net_5166), .ZN(net_5074) );
CLKBUF_X2 inst_14507 ( .A(net_13601), .Z(net_14355) );
AND2_X2 inst_9208 ( .A2(net_1908), .ZN(net_838), .A1(net_665) );
INV_X4 inst_5434 ( .ZN(net_2093), .A(net_829) );
CLKBUF_X2 inst_10418 ( .A(net_10265), .Z(net_10266) );
NAND4_X2 inst_3756 ( .A3(net_6077), .A1(net_6076), .ZN(net_4265), .A2(net_3853), .A4(net_3852) );
MUX2_X2 inst_4991 ( .A(net_9020), .Z(net_3965), .S(net_622), .B(net_609) );
CLKBUF_X2 inst_16939 ( .A(net_9409), .Z(net_16787) );
CLKBUF_X2 inst_18965 ( .A(net_12220), .Z(net_18813) );
CLKBUF_X2 inst_14993 ( .A(net_14380), .Z(net_14841) );
CLKBUF_X2 inst_16997 ( .A(net_16844), .Z(net_16845) );
CLKBUF_X2 inst_10811 ( .A(net_10658), .Z(net_10659) );
SDFF_X2 inst_1733 ( .Q(net_8144), .D(net_8144), .SI(net_2656), .SE(net_2541), .CK(net_16708) );
CLKBUF_X2 inst_9489 ( .A(net_9336), .Z(net_9337) );
AOI221_X2 inst_8832 ( .B1(net_8065), .C1(net_7861), .B2(net_6107), .ZN(net_6013), .C2(net_4400), .A(net_4297) );
CLKBUF_X2 inst_17139 ( .A(net_11069), .Z(net_16987) );
CLKBUF_X2 inst_11714 ( .A(net_11561), .Z(net_11562) );
AOI21_X2 inst_8911 ( .ZN(net_5809), .A(net_5745), .B2(net_5610), .B1(net_5258) );
NAND3_X2 inst_3900 ( .ZN(net_5638), .A1(net_5567), .A3(net_5501), .A2(net_5394) );
CLKBUF_X2 inst_18059 ( .A(net_10522), .Z(net_17907) );
SDFFR_X2 inst_2199 ( .Q(net_6483), .D(net_6483), .SE(net_2897), .SI(net_2876), .CK(net_11696), .RN(x6501) );
SDFF_X2 inst_918 ( .SI(net_8738), .Q(net_8738), .SE(net_6195), .D(net_3939), .CK(net_10502) );
NAND2_X2 inst_4751 ( .ZN(net_2716), .A2(net_1586), .A1(net_866) );
INV_X2 inst_6588 ( .A(net_6122), .ZN(net_6114) );
CLKBUF_X2 inst_16146 ( .A(net_9192), .Z(net_15994) );
CLKBUF_X2 inst_13921 ( .A(net_13768), .Z(net_13769) );
AND2_X2 inst_9177 ( .A2(net_6336), .ZN(net_5674), .A1(net_1895) );
CLKBUF_X2 inst_17846 ( .A(net_14779), .Z(net_17694) );
NAND2_X4 inst_4035 ( .ZN(net_6201), .A2(net_6090), .A1(net_6089) );
SDFF_X2 inst_1862 ( .D(net_7293), .SI(net_6950), .Q(net_6950), .SE(net_6281), .CK(net_17673) );
CLKBUF_X2 inst_14108 ( .A(net_13955), .Z(net_13956) );
CLKBUF_X2 inst_12928 ( .A(net_12775), .Z(net_12776) );
CLKBUF_X2 inst_15973 ( .A(net_10369), .Z(net_15821) );
DFFR_X1 inst_7466 ( .D(net_4403), .CK(net_9401), .RN(x6501), .Q(x1087) );
SDFFR_X2 inst_2429 ( .SE(net_2683), .D(net_1198), .SI(net_453), .Q(net_453), .CK(net_13936), .RN(x6501) );
CLKBUF_X2 inst_15292 ( .A(net_15139), .Z(net_15140) );
CLKBUF_X2 inst_18571 ( .A(net_18418), .Z(net_18419) );
CLKBUF_X2 inst_17027 ( .A(net_12823), .Z(net_16875) );
CLKBUF_X2 inst_10596 ( .A(net_10443), .Z(net_10444) );
CLKBUF_X2 inst_10463 ( .A(net_9974), .Z(net_10311) );
SDFF_X2 inst_754 ( .Q(net_8795), .D(net_8795), .SI(net_3967), .SE(net_3879), .CK(net_12253) );
CLKBUF_X2 inst_10531 ( .A(net_9989), .Z(net_10379) );
CLKBUF_X2 inst_10030 ( .A(net_9877), .Z(net_9878) );
CLKBUF_X2 inst_18696 ( .A(net_11604), .Z(net_18544) );
CLKBUF_X2 inst_18165 ( .A(net_18012), .Z(net_18013) );
CLKBUF_X2 inst_10332 ( .A(net_10179), .Z(net_10180) );
OAI22_X2 inst_2913 ( .ZN(net_4560), .A2(net_4559), .B2(net_4414), .A1(net_2522), .B1(net_301) );
AOI221_X2 inst_8783 ( .C1(net_8976), .B2(net_5538), .C2(net_5456), .ZN(net_5255), .A(net_4931), .B1(net_405) );
NOR3_X2 inst_3295 ( .ZN(net_2018), .A3(net_1698), .A2(net_1512), .A1(net_1382) );
AOI221_X2 inst_8792 ( .C1(net_7202), .C2(net_5655), .B2(net_4965), .ZN(net_4909), .A(net_4908), .B1(net_304) );
INV_X8 inst_5057 ( .ZN(net_6262), .A(net_3379) );
CLKBUF_X2 inst_16368 ( .A(net_15747), .Z(net_16216) );
AOI221_X2 inst_8828 ( .B1(net_8060), .C1(net_7856), .B2(net_6107), .ZN(net_6005), .C2(net_4400), .A(net_4303) );
DFFR_X1 inst_7394 ( .QN(net_6330), .D(net_5884), .CK(net_14229), .RN(x6501) );
CLKBUF_X2 inst_13997 ( .A(net_13844), .Z(net_13845) );
CLKBUF_X2 inst_13140 ( .A(net_12987), .Z(net_12988) );
CLKBUF_X2 inst_12998 ( .A(net_12845), .Z(net_12846) );
CLKBUF_X2 inst_16383 ( .A(net_14765), .Z(net_16231) );
OAI22_X2 inst_2923 ( .B1(net_6113), .ZN(net_2944), .B2(net_2943), .A2(net_2772), .A1(net_1429) );
AOI22_X2 inst_7957 ( .B1(net_8159), .A1(net_7717), .B2(net_6101), .A2(net_6095), .ZN(net_4170) );
SDFFR_X1 inst_2707 ( .SI(net_6811), .Q(net_6811), .SE(net_6267), .D(net_4619), .CK(net_11796), .RN(x6501) );
NAND3_X2 inst_3958 ( .A3(net_7512), .A2(net_7511), .ZN(net_2975), .A1(net_2974) );
CLKBUF_X2 inst_17543 ( .A(net_17390), .Z(net_17391) );
CLKBUF_X2 inst_10465 ( .A(net_10312), .Z(net_10313) );
CLKBUF_X2 inst_10166 ( .A(net_10013), .Z(net_10014) );
NAND2_X2 inst_4620 ( .A2(net_6144), .ZN(net_2601), .A1(net_2600) );
CLKBUF_X2 inst_12674 ( .A(net_11444), .Z(net_12522) );
CLKBUF_X2 inst_15719 ( .A(net_15566), .Z(net_15567) );
CLKBUF_X2 inst_9277 ( .A(net_9124), .Z(net_9125) );
NAND4_X2 inst_3707 ( .ZN(net_4430), .A4(net_4335), .A1(net_3720), .A2(net_3719), .A3(net_3718) );
CLKBUF_X2 inst_11869 ( .A(net_9293), .Z(net_11717) );
CLKBUF_X2 inst_14243 ( .A(net_14090), .Z(net_14091) );
CLKBUF_X2 inst_12431 ( .A(net_12278), .Z(net_12279) );
CLKBUF_X2 inst_10158 ( .A(net_10005), .Z(net_10006) );
AOI22_X2 inst_8131 ( .B1(net_8015), .A1(net_7981), .B2(net_6102), .A2(net_6097), .ZN(net_4018) );
CLKBUF_X2 inst_14767 ( .A(net_14614), .Z(net_14615) );
INV_X4 inst_5388 ( .ZN(net_1328), .A(net_1095) );
NAND2_X2 inst_4492 ( .A1(net_7204), .A2(net_5655), .ZN(net_4480) );
CLKBUF_X2 inst_13551 ( .A(net_13398), .Z(net_13399) );
CLKBUF_X2 inst_9773 ( .A(net_9620), .Z(net_9621) );
CLKBUF_X2 inst_14553 ( .A(net_14400), .Z(net_14401) );
OAI21_X2 inst_3056 ( .B2(net_8240), .B1(net_4850), .ZN(net_4751), .A(net_2605) );
CLKBUF_X2 inst_14550 ( .A(net_14397), .Z(net_14398) );
CLKBUF_X2 inst_12214 ( .A(net_12061), .Z(net_12062) );
SDFFR_X2 inst_2609 ( .Q(net_7410), .D(net_7410), .SE(net_1136), .CK(net_18653), .RN(x6501), .SI(x4919) );
SDFFR_X2 inst_2556 ( .QN(net_6351), .SE(net_2147), .D(net_2130), .SI(net_1806), .CK(net_14690), .RN(x6501) );
CLKBUF_X2 inst_15022 ( .A(net_9983), .Z(net_14870) );
INV_X4 inst_5371 ( .ZN(net_1694), .A(net_1130) );
SDFF_X2 inst_1704 ( .SI(net_7745), .Q(net_7745), .D(net_2658), .SE(net_2560), .CK(net_18843) );
NAND2_X2 inst_4604 ( .A2(net_6144), .ZN(net_2633), .A1(net_2632) );
CLKBUF_X2 inst_15156 ( .A(net_15003), .Z(net_15004) );
CLKBUF_X2 inst_15766 ( .A(net_10471), .Z(net_15614) );
XNOR2_X2 inst_161 ( .ZN(net_1847), .B(net_1846), .A(net_1752) );
CLKBUF_X2 inst_10956 ( .A(net_10803), .Z(net_10804) );
INV_X4 inst_6118 ( .A(net_7486), .ZN(net_771) );
CLKBUF_X2 inst_11287 ( .A(net_11134), .Z(net_11135) );
CLKBUF_X2 inst_9624 ( .A(net_9471), .Z(net_9472) );
CLKBUF_X2 inst_11764 ( .A(net_11611), .Z(net_11612) );
CLKBUF_X2 inst_17389 ( .A(net_13255), .Z(net_17237) );
SDFFR_X2 inst_2408 ( .SI(net_5944), .SE(net_2260), .Q(net_349), .D(net_349), .CK(net_9356), .RN(x6501) );
CLKBUF_X2 inst_10519 ( .A(net_10366), .Z(net_10367) );
CLKBUF_X2 inst_9778 ( .A(net_9207), .Z(net_9626) );
SDFF_X2 inst_1324 ( .Q(net_7812), .D(net_7812), .SE(net_2730), .SI(net_2708), .CK(net_18290) );
CLKBUF_X2 inst_15585 ( .A(net_11297), .Z(net_15433) );
CLKBUF_X2 inst_11848 ( .A(net_11695), .Z(net_11696) );
CLKBUF_X2 inst_10646 ( .A(net_10397), .Z(net_10494) );
SDFF_X2 inst_342 ( .SI(net_8593), .Q(net_8593), .SE(net_3984), .D(net_3961), .CK(net_10210) );
SDFF_X2 inst_463 ( .SI(net_8467), .Q(net_8467), .SE(net_3983), .D(net_3963), .CK(net_12350) );
CLKBUF_X2 inst_10667 ( .A(net_9299), .Z(net_10515) );
CLKBUF_X2 inst_18648 ( .A(net_9477), .Z(net_18496) );
CLKBUF_X2 inst_13571 ( .A(net_11156), .Z(net_13419) );
NAND4_X2 inst_3820 ( .ZN(net_3606), .A1(net_3407), .A2(net_3406), .A3(net_3405), .A4(net_3404) );
NAND2_X2 inst_4667 ( .ZN(net_5985), .A2(net_2328), .A1(net_2247) );
CLKBUF_X2 inst_12762 ( .A(net_11084), .Z(net_12610) );
DFFR_X2 inst_6992 ( .D(net_5898), .CK(net_11486), .RN(x6501), .Q(x2805) );
INV_X4 inst_5923 ( .A(net_6357), .ZN(net_765) );
CLKBUF_X2 inst_15857 ( .A(net_13260), .Z(net_15705) );
SDFFR_X2 inst_2158 ( .QN(net_7572), .D(net_3962), .SE(net_3144), .SI(net_582), .CK(net_13224), .RN(x6501) );
CLKBUF_X2 inst_15702 ( .A(net_11098), .Z(net_15550) );
INV_X4 inst_5560 ( .ZN(net_876), .A(net_609) );
SDFF_X2 inst_1711 ( .SI(net_7282), .Q(net_7059), .D(net_7059), .SE(net_6280), .CK(net_14909) );
CLKBUF_X2 inst_10660 ( .A(net_9107), .Z(net_10508) );
NOR2_X2 inst_3426 ( .A2(net_3093), .ZN(net_3088), .A1(net_2507) );
CLKBUF_X2 inst_16063 ( .A(net_15910), .Z(net_15911) );
CLKBUF_X2 inst_16118 ( .A(net_15965), .Z(net_15966) );
SDFF_X2 inst_2052 ( .SI(net_7779), .Q(net_7779), .D(net_2658), .SE(net_2459), .CK(net_18833) );
SDFF_X2 inst_995 ( .D(net_7334), .SI(net_6642), .Q(net_6642), .SE(net_3123), .CK(net_12033) );
AOI221_X2 inst_8850 ( .B1(net_8872), .C1(net_8317), .B2(net_6252), .C2(net_4345), .ZN(net_4342), .A(net_4255) );
CLKBUF_X2 inst_13948 ( .A(net_13795), .Z(net_13796) );
CLKBUF_X2 inst_10697 ( .A(net_10544), .Z(net_10545) );
SDFFR_X2 inst_2470 ( .D(net_6319), .SE(net_2685), .SI(net_441), .Q(net_441), .CK(net_17441), .RN(x6501) );
INV_X4 inst_6049 ( .A(net_6752), .ZN(net_498) );
NAND4_X2 inst_3857 ( .A2(net_3544), .A1(net_3309), .A4(net_3056), .A3(net_2916), .ZN(net_1435) );
CLKBUF_X2 inst_18384 ( .A(net_18231), .Z(net_18232) );
SDFF_X2 inst_1060 ( .D(net_7330), .SI(net_6638), .Q(net_6638), .SE(net_3123), .CK(net_11325) );
INV_X4 inst_5920 ( .A(net_8921), .ZN(net_2614) );
SDFF_X2 inst_900 ( .SI(net_8716), .Q(net_8716), .SE(net_6195), .D(net_3945), .CK(net_10688) );
DFFS_X1 inst_6950 ( .D(net_6145), .CK(net_13621), .SN(x6501), .Q(x801) );
CLKBUF_X2 inst_10568 ( .A(net_9686), .Z(net_10416) );
CLKBUF_X2 inst_18172 ( .A(net_18019), .Z(net_18020) );
CLKBUF_X2 inst_18123 ( .A(net_17970), .Z(net_17971) );
CLKBUF_X2 inst_14511 ( .A(net_14358), .Z(net_14359) );
MUX2_X2 inst_4949 ( .A(net_2760), .S(net_2378), .Z(net_2375), .B(net_907) );
CLKBUF_X2 inst_18835 ( .A(net_18682), .Z(net_18683) );
CLKBUF_X2 inst_19104 ( .A(net_18951), .Z(net_18952) );
CLKBUF_X2 inst_12677 ( .A(net_12524), .Z(net_12525) );
OR3_X2 inst_2807 ( .ZN(net_2848), .A2(net_2680), .A1(net_2653), .A3(net_2309) );
CLKBUF_X2 inst_13608 ( .A(net_13455), .Z(net_13456) );
INV_X4 inst_5327 ( .A(net_1812), .ZN(net_1534) );
INV_X4 inst_5423 ( .ZN(net_1127), .A(net_855) );
CLKBUF_X2 inst_9995 ( .A(net_9213), .Z(net_9843) );
AOI221_X2 inst_8803 ( .C2(net_4965), .ZN(net_4827), .A(net_4640), .B2(net_4537), .B1(net_2546), .C1(net_272) );
AOI222_X1 inst_8651 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3915), .B1(net_3011), .C1(net_3009), .A1(x13779) );
CLKBUF_X2 inst_15948 ( .A(net_12518), .Z(net_15796) );
CLKBUF_X2 inst_18683 ( .A(net_18530), .Z(net_18531) );
CLKBUF_X2 inst_10470 ( .A(net_10317), .Z(net_10318) );
AOI22_X2 inst_7882 ( .A2(net_5538), .ZN(net_4549), .B2(net_4388), .B1(net_2604), .A1(net_423) );
CLKBUF_X2 inst_11617 ( .A(net_11464), .Z(net_11465) );
CLKBUF_X2 inst_12161 ( .A(net_12008), .Z(net_12009) );
DFF_X1 inst_6767 ( .Q(net_7528), .D(net_4605), .CK(net_9542) );
AOI22_X2 inst_8084 ( .A1(net_7944), .B1(net_7774), .A2(net_6092), .B2(net_6091), .ZN(net_4061) );
SDFF_X2 inst_1225 ( .Q(net_7961), .D(net_7961), .SE(net_2755), .SI(net_2722), .CK(net_16013) );
CLKBUF_X2 inst_19029 ( .A(net_18876), .Z(net_18877) );
DFFR_X1 inst_7535 ( .Q(net_6419), .D(net_1843), .CK(net_17942), .RN(x6501) );
CLKBUF_X2 inst_12411 ( .A(net_12258), .Z(net_12259) );
CLKBUF_X2 inst_14256 ( .A(net_11677), .Z(net_14104) );
INV_X4 inst_5316 ( .ZN(net_1597), .A(net_1104) );
INV_X4 inst_5530 ( .A(net_1198), .ZN(net_660) );
CLKBUF_X2 inst_14427 ( .A(net_13864), .Z(net_14275) );
CLKBUF_X2 inst_14215 ( .A(net_14062), .Z(net_14063) );
NAND2_X2 inst_4551 ( .A1(net_3326), .ZN(net_3307), .A2(net_3305) );
CLKBUF_X2 inst_11397 ( .A(net_10393), .Z(net_11245) );
NAND2_X2 inst_4313 ( .A1(net_7056), .A2(net_5162), .ZN(net_5144) );
CLKBUF_X2 inst_13153 ( .A(net_13000), .Z(net_13001) );
NAND2_X2 inst_4714 ( .ZN(net_4369), .A1(net_1802), .A2(net_1801) );
CLKBUF_X2 inst_12898 ( .A(net_12745), .Z(net_12746) );
CLKBUF_X2 inst_16114 ( .A(net_15345), .Z(net_15962) );
OAI221_X2 inst_2956 ( .C2(net_8242), .B1(net_7585), .B2(net_4971), .C1(net_4928), .ZN(net_4912), .A(net_3240) );
NAND2_X2 inst_4713 ( .ZN(net_1804), .A1(net_1803), .A2(net_1620) );
CLKBUF_X2 inst_16071 ( .A(net_10258), .Z(net_15919) );
SDFF_X2 inst_412 ( .SI(net_8326), .Q(net_8326), .SE(net_3978), .D(net_3952), .CK(net_12908) );
INV_X4 inst_5463 ( .ZN(net_763), .A(net_762) );
CLKBUF_X2 inst_14721 ( .A(net_14568), .Z(net_14569) );
CLKBUF_X2 inst_13022 ( .A(net_12728), .Z(net_12870) );
AOI22_X2 inst_8295 ( .B1(net_8583), .A1(net_8472), .A2(net_6263), .B2(net_6262), .ZN(net_3747) );
CLKBUF_X2 inst_13969 ( .A(net_13816), .Z(net_13817) );
OAI21_X2 inst_3163 ( .B2(net_8947), .ZN(net_1726), .A(net_1725), .B1(net_1724) );
SDFFR_X2 inst_2504 ( .Q(net_8975), .D(net_8975), .SI(net_4669), .SE(net_2562), .CK(net_16629), .RN(x6501) );
CLKBUF_X2 inst_17132 ( .A(net_15883), .Z(net_16980) );
CLKBUF_X2 inst_13511 ( .A(net_12389), .Z(net_13359) );
CLKBUF_X2 inst_14076 ( .A(net_11540), .Z(net_13924) );
CLKBUF_X2 inst_14824 ( .A(net_14671), .Z(net_14672) );
CLKBUF_X2 inst_15469 ( .A(net_15316), .Z(net_15317) );
NOR2_X2 inst_3374 ( .ZN(net_5551), .A1(net_5330), .A2(net_5329) );
NAND2_X2 inst_4354 ( .A1(net_7109), .A2(net_5164), .ZN(net_5103) );
CLKBUF_X2 inst_18049 ( .A(net_17732), .Z(net_17897) );
NOR2_X2 inst_3438 ( .A2(net_3093), .ZN(net_3061), .A1(net_2929) );
CLKBUF_X2 inst_12541 ( .A(net_12388), .Z(net_12389) );
CLKBUF_X2 inst_14614 ( .A(net_12125), .Z(net_14462) );
CLKBUF_X2 inst_18781 ( .A(net_16853), .Z(net_18629) );
NAND4_X2 inst_3811 ( .ZN(net_3615), .A1(net_3443), .A2(net_3442), .A3(net_3441), .A4(net_3440) );
NAND4_X2 inst_3653 ( .A4(net_6034), .A1(net_6033), .ZN(net_4612), .A2(net_4174), .A3(net_4173) );
CLKBUF_X2 inst_18694 ( .A(net_18541), .Z(net_18542) );
DFFS_X1 inst_6959 ( .D(net_2586), .CK(net_16572), .SN(x6501), .Q(x677) );
CLKBUF_X2 inst_15652 ( .A(net_15499), .Z(net_15500) );
AOI22_X2 inst_8213 ( .B1(net_8572), .A1(net_8461), .A2(net_6263), .B2(net_6262), .ZN(net_3823) );
CLKBUF_X2 inst_10700 ( .A(net_10547), .Z(net_10548) );
CLKBUF_X2 inst_16187 ( .A(net_16034), .Z(net_16035) );
CLKBUF_X2 inst_15438 ( .A(net_15285), .Z(net_15286) );
SDFF_X2 inst_1241 ( .Q(net_7968), .D(net_7968), .SE(net_2755), .SI(net_2710), .CK(net_14191) );
SDFF_X2 inst_1038 ( .SI(net_7316), .Q(net_6690), .D(net_6690), .SE(net_3125), .CK(net_9863) );
CLKBUF_X2 inst_15418 ( .A(net_13234), .Z(net_15266) );
SDFF_X2 inst_940 ( .SI(net_7320), .Q(net_6661), .D(net_6661), .SE(net_3126), .CK(net_12146) );
CLKBUF_X2 inst_9417 ( .A(net_9062), .Z(net_9265) );
CLKBUF_X2 inst_11705 ( .A(net_9235), .Z(net_11553) );
CLKBUF_X2 inst_11641 ( .A(net_11488), .Z(net_11489) );
NOR2_X2 inst_3595 ( .A1(net_7522), .A2(net_1501), .ZN(net_892) );
CLKBUF_X2 inst_11830 ( .A(net_11677), .Z(net_11678) );
NAND2_X2 inst_4876 ( .A2(net_3274), .ZN(net_1065), .A1(net_544) );
AOI22_X2 inst_8103 ( .B2(net_8110), .A1(net_7770), .B1(net_6108), .A2(net_6096), .ZN(net_4045) );
CLKBUF_X1 inst_7732 ( .A(x192486), .Z(x1062) );
AOI211_X2 inst_9008 ( .C2(net_5538), .ZN(net_5458), .B(net_4977), .A(net_4976), .C1(net_762) );
NAND2_X2 inst_4362 ( .A1(net_7151), .A2(net_5166), .ZN(net_5095) );
CLKBUF_X2 inst_9581 ( .A(net_9428), .Z(net_9429) );
CLKBUF_X2 inst_15761 ( .A(net_15321), .Z(net_15609) );
CLKBUF_X2 inst_12608 ( .A(net_11914), .Z(net_12456) );
NAND2_X2 inst_4369 ( .A1(net_7113), .A2(net_5164), .ZN(net_5088) );
CLKBUF_X2 inst_17869 ( .A(net_15748), .Z(net_17717) );
CLKBUF_X2 inst_11899 ( .A(net_11224), .Z(net_11747) );
CLKBUF_X2 inst_11236 ( .A(net_11083), .Z(net_11084) );
CLKBUF_X2 inst_13076 ( .A(net_12642), .Z(net_12924) );
NAND3_X2 inst_4007 ( .A3(net_7348), .ZN(net_1475), .A2(net_1085), .A1(net_1060) );
SDFF_X2 inst_879 ( .Q(net_8591), .D(net_8591), .SI(net_3949), .SE(net_3878), .CK(net_12779) );
CLKBUF_X2 inst_17325 ( .A(net_10201), .Z(net_17173) );
CLKBUF_X2 inst_17105 ( .A(net_12152), .Z(net_16953) );
NAND2_X2 inst_4291 ( .A1(net_7080), .ZN(net_5169), .A2(net_5164) );
INV_X4 inst_5692 ( .ZN(net_2641), .A(net_156) );
CLKBUF_X2 inst_17603 ( .A(net_14521), .Z(net_17451) );
SDFF_X2 inst_629 ( .SI(net_8542), .Q(net_8542), .SE(net_3979), .D(net_3942), .CK(net_12795) );
NAND2_X2 inst_4903 ( .A2(net_7387), .ZN(net_616), .A1(net_176) );
SDFF_X2 inst_1100 ( .D(net_7330), .SI(net_6539), .Q(net_6539), .SE(net_3086), .CK(net_11321) );
CLKBUF_X2 inst_10872 ( .A(net_10358), .Z(net_10720) );
CLKBUF_X2 inst_18037 ( .A(net_15066), .Z(net_17885) );
CLKBUF_X2 inst_15105 ( .A(net_14491), .Z(net_14953) );
CLKBUF_X2 inst_18372 ( .A(net_18219), .Z(net_18220) );
NOR2_X2 inst_3383 ( .ZN(net_5542), .A1(net_5293), .A2(net_5292) );
CLKBUF_X2 inst_15682 ( .A(net_15529), .Z(net_15530) );
SDFF_X2 inst_1191 ( .D(net_7311), .SI(net_6553), .Q(net_6553), .SE(net_3070), .CK(net_9890) );
CLKBUF_X2 inst_18307 ( .A(net_18154), .Z(net_18155) );
SDFF_X2 inst_533 ( .Q(net_8858), .D(net_8858), .SI(net_3947), .SE(net_3936), .CK(net_12455) );
SDFFR_X2 inst_2478 ( .Q(net_8989), .D(net_8989), .SI(net_2608), .SE(net_2562), .CK(net_16644), .RN(x6501) );
MUX2_X2 inst_4972 ( .S(net_6325), .Z(net_4956), .A(net_592), .B(x4932) );
SDFFR_X1 inst_2751 ( .SI(net_9025), .Q(net_9025), .D(net_7454), .SE(net_3208), .CK(net_12928), .RN(x6501) );
CLKBUF_X2 inst_16928 ( .A(net_15571), .Z(net_16776) );
SDFF_X2 inst_1760 ( .SI(net_7761), .Q(net_7761), .D(net_2749), .SE(net_2560), .CK(net_13749) );
SDFF_X2 inst_1874 ( .D(net_7277), .SI(net_6974), .Q(net_6974), .SE(net_6283), .CK(net_14613) );
SDFF_X2 inst_2022 ( .SI(net_7930), .Q(net_7930), .D(net_2712), .SE(net_2461), .CK(net_17111) );
NAND3_X2 inst_3960 ( .A1(net_6201), .A3(net_6170), .A2(net_6093), .ZN(net_6088) );
OR2_X4 inst_2821 ( .ZN(net_4950), .A1(net_4385), .A2(net_4318) );
SDFF_X2 inst_1095 ( .D(net_7311), .SI(net_6520), .Q(net_6520), .SE(net_3086), .CK(net_9925) );
AOI22_X2 inst_8042 ( .B1(net_8204), .A1(net_7694), .B2(net_6099), .A2(net_4399), .ZN(net_4097) );
CLKBUF_X2 inst_16738 ( .A(net_16585), .Z(net_16586) );
CLKBUF_X2 inst_10516 ( .A(net_9318), .Z(net_10364) );
CLKBUF_X2 inst_10096 ( .A(net_9203), .Z(net_9944) );
AND2_X4 inst_9052 ( .ZN(net_3360), .A2(net_3356), .A1(net_3328) );
SDFFR_X2 inst_2439 ( .D(net_4457), .SE(net_2313), .SI(net_421), .Q(net_421), .CK(net_17281), .RN(x6501) );
XNOR2_X2 inst_176 ( .ZN(net_1758), .B(net_1757), .A(net_1445) );
OR2_X4 inst_2826 ( .ZN(net_3572), .A1(net_3570), .A2(net_3529) );
AND2_X4 inst_9069 ( .ZN(net_3520), .A1(net_3250), .A2(net_3216) );
CLKBUF_X2 inst_10894 ( .A(net_9076), .Z(net_10742) );
SDFF_X2 inst_1336 ( .SI(net_7680), .Q(net_7680), .SE(net_2714), .D(net_2584), .CK(net_15616) );
INV_X4 inst_5472 ( .ZN(net_1151), .A(net_1074) );
CLKBUF_X2 inst_10387 ( .A(net_10234), .Z(net_10235) );
SDFF_X2 inst_1665 ( .SI(net_7760), .Q(net_7760), .D(net_2712), .SE(net_2560), .CK(net_13767) );
NAND2_X2 inst_4500 ( .ZN(net_4414), .A2(net_4397), .A1(net_4383) );
CLKBUF_X2 inst_13962 ( .A(net_13809), .Z(net_13810) );
NAND2_X2 inst_4763 ( .A1(net_6117), .ZN(net_1706), .A2(net_1705) );
CLKBUF_X2 inst_17224 ( .A(net_17071), .Z(net_17072) );
SDFF_X2 inst_780 ( .SI(net_8349), .Q(net_8349), .D(net_3973), .SE(net_3880), .CK(net_10827) );
INV_X4 inst_5626 ( .A(net_7666), .ZN(net_917) );
DFF_X1 inst_6783 ( .Q(net_7532), .D(net_4587), .CK(net_11963) );
AOI22_X2 inst_8255 ( .A1(net_8614), .B1(net_8429), .A2(net_3864), .B2(net_3863), .ZN(net_3783) );
CLKBUF_X2 inst_12016 ( .A(net_11863), .Z(net_11864) );
NAND3_X2 inst_3967 ( .ZN(net_2734), .A1(net_2315), .A3(net_2314), .A2(net_1885) );
CLKBUF_X2 inst_19099 ( .A(net_10261), .Z(net_18947) );
CLKBUF_X2 inst_16769 ( .A(net_16616), .Z(net_16617) );
AOI221_X4 inst_8722 ( .B1(net_8723), .C1(net_8501), .B2(net_4350), .C2(net_4349), .ZN(net_4344), .A(net_4257) );
NAND4_X2 inst_3669 ( .A4(net_6024), .A1(net_6023), .ZN(net_4596), .A2(net_4078), .A3(net_4077) );
SDFF_X2 inst_1767 ( .D(net_7287), .SI(net_6864), .Q(net_6864), .SE(net_6282), .CK(net_14901) );
CLKBUF_X2 inst_13564 ( .A(net_9850), .Z(net_13412) );
CLKBUF_X2 inst_16087 ( .A(net_15934), .Z(net_15935) );
SDFFR_X2 inst_2361 ( .SE(net_2260), .Q(net_337), .D(net_337), .CK(net_9308), .RN(x6501), .SI(x2308) );
CLKBUF_X2 inst_11497 ( .A(net_11344), .Z(net_11345) );
CLKBUF_X2 inst_10237 ( .A(net_10084), .Z(net_10085) );
INV_X4 inst_6006 ( .A(net_6352), .ZN(net_512) );
CLKBUF_X2 inst_14652 ( .A(net_14499), .Z(net_14500) );
DFF_X1 inst_6802 ( .QN(net_8248), .D(net_4431), .CK(net_16272) );
CLKBUF_X2 inst_16797 ( .A(net_13781), .Z(net_16645) );
SDFF_X2 inst_694 ( .Q(net_8853), .D(net_8853), .SI(net_3943), .SE(net_3936), .CK(net_13339) );
CLKBUF_X2 inst_17025 ( .A(net_12352), .Z(net_16873) );
CLKBUF_X2 inst_15689 ( .A(net_15536), .Z(net_15537) );
INV_X4 inst_5574 ( .A(net_7605), .ZN(net_1930) );
INV_X2 inst_6382 ( .A(net_1694), .ZN(net_1471) );
SDFFR_X2 inst_2498 ( .Q(net_8974), .D(net_8974), .SI(net_2624), .SE(net_2562), .CK(net_14794), .RN(x6501) );
CLKBUF_X2 inst_17274 ( .A(net_15446), .Z(net_17122) );
CLKBUF_X2 inst_12402 ( .A(net_12249), .Z(net_12250) );
OAI21_X2 inst_3154 ( .B2(net_1984), .ZN(net_1980), .A(net_1979), .B1(net_752) );
INV_X4 inst_5396 ( .A(net_1661), .ZN(net_914) );
CLKBUF_X2 inst_9394 ( .A(net_9186), .Z(net_9242) );
CLKBUF_X2 inst_15531 ( .A(net_11101), .Z(net_15379) );
AOI22_X2 inst_7814 ( .A2(net_8247), .B2(net_6144), .A1(net_4764), .ZN(net_4744), .B1(net_4743) );
CLKBUF_X2 inst_17390 ( .A(net_17237), .Z(net_17238) );
CLKBUF_X2 inst_16767 ( .A(net_16614), .Z(net_16615) );
CLKBUF_X2 inst_16271 ( .A(net_14734), .Z(net_16119) );
CLKBUF_X2 inst_12071 ( .A(net_11557), .Z(net_11919) );
SDFF_X2 inst_787 ( .SI(net_8357), .Q(net_8357), .D(net_3942), .SE(net_3880), .CK(net_12587) );
NAND2_X2 inst_4396 ( .A1(net_7085), .A2(net_5164), .ZN(net_5061) );
CLKBUF_X2 inst_11211 ( .A(net_10898), .Z(net_11059) );
CLKBUF_X2 inst_12958 ( .A(net_9496), .Z(net_12806) );
CLKBUF_X2 inst_18214 ( .A(net_18061), .Z(net_18062) );
CLKBUF_X2 inst_15541 ( .A(net_15388), .Z(net_15389) );
CLKBUF_X2 inst_14439 ( .A(net_9853), .Z(net_14287) );
SDFF_X2 inst_825 ( .SI(net_8518), .Q(net_8518), .D(net_3948), .SE(net_3884), .CK(net_13391) );
SDFFR_X2 inst_2586 ( .D(net_7392), .QN(net_7252), .SI(net_1951), .SE(net_1379), .CK(net_18317), .RN(x6501) );
AOI22_X2 inst_7928 ( .B1(net_7908), .A1(net_7806), .B2(net_6103), .A2(net_4398), .ZN(net_4196) );
CLKBUF_X2 inst_17684 ( .A(net_14892), .Z(net_17532) );
CLKBUF_X2 inst_15310 ( .A(net_15157), .Z(net_15158) );
CLKBUF_X2 inst_12886 ( .A(net_12733), .Z(net_12734) );
SDFF_X2 inst_1892 ( .D(net_7291), .SI(net_6868), .Q(net_6868), .SE(net_6282), .CK(net_17665) );
AOI22_X2 inst_7860 ( .B2(net_4881), .A2(net_4809), .ZN(net_4581), .A1(net_343), .B1(net_249) );
CLKBUF_X2 inst_11404 ( .A(net_10014), .Z(net_11252) );
SDFF_X2 inst_726 ( .SI(net_8498), .Q(net_8498), .D(net_3944), .SE(net_3884), .CK(net_13103) );
CLKBUF_X2 inst_18112 ( .A(net_12959), .Z(net_17960) );
CLKBUF_X2 inst_18436 ( .A(net_12753), .Z(net_18284) );
CLKBUF_X2 inst_10583 ( .A(net_10430), .Z(net_10431) );
CLKBUF_X2 inst_18988 ( .A(net_18835), .Z(net_18836) );
NAND2_X2 inst_4726 ( .A1(net_7367), .ZN(net_2056), .A2(net_1782) );
AOI22_X2 inst_8073 ( .B1(net_8141), .A1(net_7903), .A2(net_6098), .B2(net_4190), .ZN(net_4071) );
CLKBUF_X2 inst_18623 ( .A(net_18470), .Z(net_18471) );
XNOR2_X2 inst_320 ( .B(net_7390), .ZN(net_941), .A(net_571) );
CLKBUF_X2 inst_16861 ( .A(net_12498), .Z(net_16709) );
XOR2_X2 inst_1 ( .B(net_3388), .Z(net_3238), .A(net_3096) );
CLKBUF_X2 inst_16327 ( .A(net_12985), .Z(net_16175) );
SDFF_X2 inst_1891 ( .D(net_7274), .SI(net_7011), .Q(net_7011), .SE(net_6277), .CK(net_14093) );
CLKBUF_X2 inst_12794 ( .A(net_12641), .Z(net_12642) );
NAND2_X2 inst_4558 ( .A1(net_6387), .A2(net_6184), .ZN(net_3252) );
CLKBUF_X2 inst_14862 ( .A(net_11009), .Z(net_14710) );
CLKBUF_X2 inst_14525 ( .A(net_10866), .Z(net_14373) );
CLKBUF_X2 inst_19175 ( .A(net_19022), .Z(net_19023) );
CLKBUF_X2 inst_17411 ( .A(net_16862), .Z(net_17259) );
OAI21_X2 inst_3063 ( .B2(net_8249), .B1(net_4850), .ZN(net_4741), .A(net_2621) );
CLKBUF_X2 inst_13881 ( .A(net_13255), .Z(net_13729) );
CLKBUF_X2 inst_17770 ( .A(net_9207), .Z(net_17618) );
CLKBUF_X2 inst_17691 ( .A(net_17538), .Z(net_17539) );
SDFF_X2 inst_1812 ( .D(net_7302), .SI(net_7039), .Q(net_7039), .SE(net_6277), .CK(net_15421) );
CLKBUF_X2 inst_15036 ( .A(net_14883), .Z(net_14884) );
CLKBUF_X2 inst_14608 ( .A(net_14455), .Z(net_14456) );
CLKBUF_X2 inst_17258 ( .A(net_17105), .Z(net_17106) );
CLKBUF_X2 inst_12726 ( .A(net_9797), .Z(net_12574) );
CLKBUF_X2 inst_13066 ( .A(net_12913), .Z(net_12914) );
NAND2_X2 inst_4721 ( .A1(net_7369), .ZN(net_1985), .A2(net_1783) );
CLKBUF_X2 inst_13601 ( .A(net_9404), .Z(net_13449) );
INV_X16 inst_6638 ( .ZN(net_3935), .A(net_3350) );
CLKBUF_X2 inst_13019 ( .A(net_12866), .Z(net_12867) );
SDFFR_X2 inst_2207 ( .D(net_2483), .SE(net_2476), .SI(net_386), .Q(net_386), .CK(net_11576), .RN(x6501) );
AOI22_X2 inst_7841 ( .A2(net_5595), .ZN(net_4668), .B2(net_4388), .B1(net_2622), .A1(net_311) );
CLKBUF_X2 inst_16254 ( .A(net_12143), .Z(net_16102) );
CLKBUF_X2 inst_10088 ( .A(net_9935), .Z(net_9936) );
CLKBUF_X2 inst_17086 ( .A(net_9063), .Z(net_16934) );
CLKBUF_X2 inst_15692 ( .A(net_15539), .Z(net_15540) );
INV_X4 inst_5902 ( .A(net_6377), .ZN(net_532) );
DFFR_X2 inst_7322 ( .D(net_6415), .Q(net_6406), .CK(net_11925), .RN(x6501) );
NAND3_X2 inst_3892 ( .ZN(net_5646), .A1(net_5575), .A3(net_5509), .A2(net_5426) );
CLKBUF_X2 inst_16265 ( .A(net_16112), .Z(net_16113) );
CLKBUF_X2 inst_14906 ( .A(net_11628), .Z(net_14754) );
AOI221_X2 inst_8829 ( .C1(net_8164), .B1(net_7722), .C2(net_6101), .B2(net_6095), .ZN(net_6007), .A(net_4301) );
NAND3_X2 inst_3930 ( .ZN(net_5585), .A1(net_5458), .A2(net_4691), .A3(net_4661) );
OR2_X2 inst_2867 ( .ZN(net_5876), .A1(net_2413), .A2(net_257) );
CLKBUF_X2 inst_16388 ( .A(net_9205), .Z(net_16236) );
CLKBUF_X2 inst_9768 ( .A(net_9615), .Z(net_9616) );
AOI22_X2 inst_7953 ( .B1(net_7921), .A1(net_7819), .B2(net_6103), .A2(net_4398), .ZN(net_4174) );
CLKBUF_X2 inst_17147 ( .A(net_16994), .Z(net_16995) );
CLKBUF_X2 inst_14235 ( .A(net_13974), .Z(net_14083) );
NOR3_X2 inst_3305 ( .ZN(net_2046), .A3(net_1521), .A2(net_1347), .A1(net_751) );
CLKBUF_X2 inst_14637 ( .A(net_14484), .Z(net_14485) );
CLKBUF_X2 inst_10153 ( .A(net_9352), .Z(net_10001) );
SDFF_X2 inst_710 ( .SI(net_8666), .Q(net_8666), .D(net_3948), .SE(net_3885), .CK(net_13470) );
SDFF_X2 inst_941 ( .SI(net_7321), .Q(net_6695), .D(net_6695), .SE(net_3125), .CK(net_12142) );
NOR2_X2 inst_3350 ( .ZN(net_5575), .A1(net_5428), .A2(net_5427) );
AOI22_X2 inst_8398 ( .B1(net_8785), .A1(net_8526), .A2(net_3861), .B2(net_3860), .ZN(net_3654) );
XOR2_X2 inst_56 ( .A(net_3921), .Z(net_974), .B(net_511) );
DFF_X1 inst_6835 ( .Q(net_6427), .D(net_3613), .CK(net_17981) );
XNOR2_X2 inst_308 ( .B(net_8289), .ZN(net_963), .A(net_958) );
SDFF_X2 inst_1546 ( .Q(net_8002), .D(net_8002), .SI(net_2710), .SE(net_2542), .CK(net_16502) );
DFFR_X2 inst_7208 ( .D(net_2368), .QN(net_213), .CK(net_17884), .RN(x6501) );
CLKBUF_X2 inst_11224 ( .A(net_9894), .Z(net_11072) );
SDFF_X2 inst_455 ( .SI(net_8457), .Q(net_8457), .SE(net_3983), .D(net_3945), .CK(net_11106) );
AOI22_X2 inst_8449 ( .B1(net_6669), .A1(net_6636), .A2(net_6213), .B2(net_6138), .ZN(net_3491) );
CLKBUF_X2 inst_10015 ( .A(net_9862), .Z(net_9863) );
SDFF_X2 inst_1694 ( .SI(net_7294), .Q(net_7071), .D(net_7071), .SE(net_6280), .CK(net_17693) );
CLKBUF_X2 inst_17153 ( .A(net_17000), .Z(net_17001) );
CLKBUF_X2 inst_17158 ( .A(net_17005), .Z(net_17006) );
SDFFR_X2 inst_2540 ( .QN(net_6363), .SE(net_2147), .SI(net_1945), .D(net_695), .CK(net_14759), .RN(x6501) );
DFF_X1 inst_6833 ( .Q(net_6453), .D(net_3615), .CK(net_15159) );
CLKBUF_X2 inst_13298 ( .A(net_13145), .Z(net_13146) );
CLKBUF_X2 inst_17231 ( .A(net_17078), .Z(net_17079) );
DFFR_X2 inst_7052 ( .QN(net_7502), .D(net_4830), .CK(net_16676), .RN(x6501) );
INV_X2 inst_6602 ( .A(net_6160), .ZN(net_6159) );
AOI22_X2 inst_8114 ( .B1(net_8115), .A1(net_7877), .A2(net_6098), .B2(net_4190), .ZN(net_4034) );
OAI21_X2 inst_3024 ( .ZN(net_4972), .B2(net_4971), .A(net_4767), .B1(net_750) );
CLKBUF_X2 inst_18406 ( .A(net_18253), .Z(net_18254) );
AOI22_X2 inst_8454 ( .B1(net_6670), .A1(net_6637), .A2(net_6213), .B2(net_6138), .ZN(net_3486) );
CLKBUF_X2 inst_17942 ( .A(net_17789), .Z(net_17790) );
CLKBUF_X2 inst_11860 ( .A(net_11707), .Z(net_11708) );
CLKBUF_X2 inst_16370 ( .A(net_16217), .Z(net_16218) );
NAND3_X2 inst_3951 ( .ZN(net_3364), .A2(net_3363), .A3(net_3362), .A1(net_1378) );
AOI22_X2 inst_8240 ( .B1(net_8779), .A1(net_8520), .A2(net_3861), .B2(net_3860), .ZN(net_3797) );
CLKBUF_X2 inst_16337 ( .A(net_16184), .Z(net_16185) );
NAND2_X2 inst_4282 ( .A1(net_7006), .A2(net_5249), .ZN(net_5178) );
INV_X4 inst_5428 ( .A(net_8217), .ZN(net_1130) );
CLKBUF_X2 inst_18197 ( .A(net_18044), .Z(net_18045) );
OAI22_X2 inst_2943 ( .A1(net_2043), .ZN(net_1875), .A2(net_1788), .B1(net_1684), .B2(net_1136) );
SDFF_X2 inst_1593 ( .Q(net_8124), .D(net_8124), .SI(net_2574), .SE(net_2541), .CK(net_18378) );
CLKBUF_X2 inst_18595 ( .A(net_11762), .Z(net_18443) );
SDFF_X2 inst_724 ( .SI(net_8512), .Q(net_8512), .D(net_3940), .SE(net_3884), .CK(net_13468) );
CLKBUF_X2 inst_17526 ( .A(net_17373), .Z(net_17374) );
CLKBUF_X2 inst_14869 ( .A(net_14716), .Z(net_14717) );
SDFF_X2 inst_975 ( .SI(net_7339), .Q(net_6746), .D(net_6746), .SE(net_3124), .CK(net_11913) );
CLKBUF_X2 inst_15546 ( .A(net_15393), .Z(net_15394) );
CLKBUF_X2 inst_16677 ( .A(net_16524), .Z(net_16525) );
CLKBUF_X2 inst_13683 ( .A(net_10536), .Z(net_13531) );
OAI211_X2 inst_3191 ( .C2(net_8890), .ZN(net_3902), .B(net_3901), .C1(net_3587), .A(net_1407) );
SDFFR_X1 inst_2789 ( .D(net_7392), .Q(net_7289), .SI(net_1951), .SE(net_1327), .CK(net_15363), .RN(x6501) );
AOI22_X2 inst_7792 ( .A2(net_6187), .B2(net_5463), .ZN(net_4806), .B1(net_441), .A1(net_204) );
CLKBUF_X2 inst_9504 ( .A(net_9351), .Z(net_9352) );
INV_X4 inst_5714 ( .A(net_7598), .ZN(net_1004) );
CLKBUF_X2 inst_10110 ( .A(net_9957), .Z(net_9958) );
CLKBUF_X2 inst_10783 ( .A(net_10630), .Z(net_10631) );
SDFF_X2 inst_1804 ( .D(net_7264), .SI(net_7001), .Q(net_7001), .SE(net_6277), .CK(net_14155) );
INV_X2 inst_6418 ( .ZN(net_781), .A(net_780) );
CLKBUF_X2 inst_18778 ( .A(net_18625), .Z(net_18626) );
CLKBUF_X2 inst_11037 ( .A(net_10884), .Z(net_10885) );
SDFFR_X2 inst_2183 ( .QN(net_7521), .SE(net_2910), .SI(net_2909), .D(net_1076), .CK(net_9616), .RN(x6501) );
CLKBUF_X2 inst_11981 ( .A(net_9147), .Z(net_11829) );
INV_X4 inst_5068 ( .ZN(net_5877), .A(net_5839) );
SDFFR_X1 inst_2659 ( .D(net_6781), .SE(net_4506), .CK(net_11413), .RN(x6501), .SI(x1428), .Q(x1428) );
INV_X2 inst_6545 ( .A(net_7364), .ZN(net_2242) );
CLKBUF_X2 inst_13878 ( .A(net_13118), .Z(net_13726) );
INV_X8 inst_5018 ( .ZN(net_5609), .A(net_4379) );
CLKBUF_X2 inst_11609 ( .A(net_10203), .Z(net_11457) );
CLKBUF_X2 inst_18144 ( .A(net_17991), .Z(net_17992) );
INV_X4 inst_5641 ( .A(net_7614), .ZN(net_2807) );
CLKBUF_X2 inst_11134 ( .A(net_9405), .Z(net_10982) );
CLKBUF_X2 inst_18708 ( .A(net_18555), .Z(net_18556) );
CLKBUF_X2 inst_18814 ( .A(net_13582), .Z(net_18662) );
SDFF_X2 inst_1155 ( .SI(net_7337), .Q(net_6612), .D(net_6612), .SE(net_3069), .CK(net_9448) );
XNOR2_X2 inst_207 ( .ZN(net_1493), .B(net_1492), .A(net_1346) );
CLKBUF_X2 inst_16169 ( .A(net_14733), .Z(net_16017) );
AOI21_X2 inst_8886 ( .B2(net_5871), .ZN(net_5812), .A(net_5807), .B1(x420) );
CLKBUF_X2 inst_14467 ( .A(net_11497), .Z(net_14315) );
CLKBUF_X2 inst_18096 ( .A(net_15086), .Z(net_17944) );
CLKBUF_X2 inst_10490 ( .A(net_10337), .Z(net_10338) );
CLKBUF_X2 inst_9615 ( .A(net_9462), .Z(net_9463) );
CLKBUF_X2 inst_9912 ( .A(net_9759), .Z(net_9760) );
SDFF_X2 inst_1215 ( .Q(net_7969), .D(net_7969), .SE(net_2755), .SI(net_2639), .CK(net_16882) );
CLKBUF_X2 inst_9303 ( .A(net_9071), .Z(net_9151) );
XNOR2_X2 inst_131 ( .ZN(net_2816), .B(net_2754), .A(net_2753) );
CLKBUF_X2 inst_15353 ( .A(net_15200), .Z(net_15201) );
INV_X4 inst_6104 ( .A(net_7379), .ZN(net_1745) );
CLKBUF_X2 inst_16412 ( .A(net_16259), .Z(net_16260) );
XOR2_X2 inst_47 ( .A(net_3129), .Z(net_1017), .B(net_1016) );
CLKBUF_X2 inst_12360 ( .A(net_12207), .Z(net_12208) );
CLKBUF_X2 inst_14958 ( .A(net_14805), .Z(net_14806) );
SDFF_X2 inst_1984 ( .SI(net_6876), .Q(net_6876), .SE(net_6282), .D(net_2544), .CK(net_15865) );
INV_X4 inst_5231 ( .ZN(net_5745), .A(net_2252) );
CLKBUF_X2 inst_14567 ( .A(net_13047), .Z(net_14415) );
CLKBUF_X2 inst_9458 ( .A(net_9101), .Z(net_9306) );
CLKBUF_X2 inst_15563 ( .A(net_15410), .Z(net_15411) );
INV_X2 inst_6520 ( .ZN(net_787), .A(net_220) );
CLKBUF_X2 inst_14356 ( .A(net_11314), .Z(net_14204) );
CLKBUF_X2 inst_12397 ( .A(net_12244), .Z(net_12245) );
NAND2_X2 inst_4101 ( .ZN(net_5432), .A1(net_5155), .A2(net_5154) );
CLKBUF_X2 inst_10316 ( .A(net_10163), .Z(net_10164) );
CLKBUF_X2 inst_9469 ( .A(net_9316), .Z(net_9317) );
NAND2_X2 inst_4792 ( .ZN(net_1992), .A1(net_1129), .A2(net_716) );
CLKBUF_X2 inst_14027 ( .A(net_10360), .Z(net_13875) );
CLKBUF_X2 inst_18249 ( .A(net_16785), .Z(net_18097) );
CLKBUF_X2 inst_17078 ( .A(net_16925), .Z(net_16926) );
CLKBUF_X2 inst_12738 ( .A(net_12585), .Z(net_12586) );
SDFF_X2 inst_434 ( .Q(net_8762), .D(net_8762), .SE(net_3982), .SI(net_3956), .CK(net_13283) );
NOR2_X2 inst_3455 ( .A1(net_3023), .ZN(net_2877), .A2(net_2816) );
CLKBUF_X2 inst_14099 ( .A(net_13946), .Z(net_13947) );
SDFF_X2 inst_1392 ( .SI(net_7277), .Q(net_7094), .D(net_7094), .SE(net_6278), .CK(net_17399) );
DFFR_X1 inst_7376 ( .D(net_5908), .CK(net_16786), .RN(x6501), .Q(x508) );
CLKBUF_X2 inst_11816 ( .A(net_11663), .Z(net_11664) );
NAND2_X4 inst_4044 ( .ZN(net_2560), .A1(net_2269), .A2(net_2268) );
CLKBUF_X2 inst_18926 ( .A(net_18773), .Z(net_18774) );
CLKBUF_X2 inst_17116 ( .A(net_11118), .Z(net_16964) );
CLKBUF_X2 inst_16971 ( .A(net_16818), .Z(net_16819) );
CLKBUF_X2 inst_16282 ( .A(net_11650), .Z(net_16130) );
CLKBUF_X2 inst_16697 ( .A(net_16544), .Z(net_16545) );
SDFF_X2 inst_1476 ( .SI(net_7271), .Q(net_7128), .D(net_7128), .SE(net_6279), .CK(net_16840) );
AOI22_X2 inst_8265 ( .B1(net_8764), .A1(net_8394), .A2(net_3867), .B2(net_3866), .ZN(net_3773) );
SDFFR_X2 inst_2249 ( .D(net_7378), .SE(net_2802), .SI(net_187), .Q(net_187), .CK(net_14988), .RN(x6501) );
CLKBUF_X2 inst_18187 ( .A(net_16896), .Z(net_18035) );
CLKBUF_X2 inst_13773 ( .A(net_13620), .Z(net_13621) );
AOI21_X2 inst_8995 ( .B2(net_1650), .ZN(net_1433), .A(net_1032), .B1(net_201) );
INV_X4 inst_5404 ( .ZN(net_1098), .A(net_878) );
SDFFR_X2 inst_2390 ( .SE(net_2260), .Q(net_382), .D(net_382), .CK(net_9360), .RN(x6501), .SI(x1244) );
CLKBUF_X2 inst_17315 ( .A(net_17162), .Z(net_17163) );
INV_X4 inst_6033 ( .A(net_7344), .ZN(net_703) );
CLKBUF_X2 inst_17592 ( .A(net_12322), .Z(net_17440) );
CLKBUF_X2 inst_15149 ( .A(net_14996), .Z(net_14997) );
CLKBUF_X2 inst_14305 ( .A(net_9300), .Z(net_14153) );
AOI22_X2 inst_8424 ( .B1(net_6530), .A1(net_6497), .A2(net_6137), .B2(net_6104), .ZN(net_3517) );
NAND3_X4 inst_3871 ( .A1(net_6261), .A3(net_6190), .ZN(net_4709), .A2(net_4708) );
CLKBUF_X2 inst_9268 ( .A(net_9115), .Z(net_9116) );
NAND2_X2 inst_4449 ( .A1(net_6849), .A2(net_5016), .ZN(net_4978) );
INV_X4 inst_6077 ( .A(net_6363), .ZN(net_695) );
SDFF_X2 inst_2045 ( .SI(net_7929), .Q(net_7929), .D(net_2713), .SE(net_2461), .CK(net_14377) );
CLKBUF_X2 inst_17807 ( .A(net_17654), .Z(net_17655) );
CLKBUF_X2 inst_11746 ( .A(net_10240), .Z(net_11594) );
SDFF_X2 inst_1311 ( .Q(net_8088), .D(net_8088), .SE(net_2707), .SI(net_2584), .CK(net_18885) );
CLKBUF_X2 inst_9307 ( .A(net_9154), .Z(net_9155) );
DFFR_X2 inst_7185 ( .QN(net_8959), .D(net_2490), .CK(net_15072), .RN(x6501) );
NOR2_X2 inst_3415 ( .ZN(net_3305), .A2(net_3175), .A1(net_1110) );
CLKBUF_X2 inst_9534 ( .A(net_9381), .Z(net_9382) );
CLKBUF_X2 inst_16667 ( .A(net_16514), .Z(net_16515) );
CLKBUF_X2 inst_10780 ( .A(net_10627), .Z(net_10628) );
NAND2_X2 inst_4654 ( .A1(net_2555), .ZN(net_2323), .A2(net_2220) );
SDFF_X2 inst_1640 ( .SI(net_7704), .Q(net_7704), .D(net_2721), .SE(net_2559), .CK(net_15756) );
CLKBUF_X2 inst_11359 ( .A(net_11206), .Z(net_11207) );
CLKBUF_X2 inst_13928 ( .A(net_13775), .Z(net_13776) );
CLKBUF_X2 inst_15127 ( .A(net_13489), .Z(net_14975) );
NAND2_X2 inst_4747 ( .ZN(net_2639), .A1(net_1780), .A2(net_1586) );
DFFR_X1 inst_7571 ( .Q(net_7619), .D(net_7616), .CK(net_11183), .RN(x6501) );
NAND2_X2 inst_4630 ( .A2(net_5871), .ZN(net_2515), .A1(x626) );
SDFFR_X2 inst_2509 ( .Q(net_8995), .D(net_8995), .SI(net_2596), .SE(net_2562), .CK(net_14527), .RN(x6501) );
INV_X4 inst_5971 ( .A(net_8897), .ZN(net_1150) );
OAI21_X2 inst_3091 ( .B2(net_2897), .ZN(net_2895), .A(net_2894), .B1(net_1145) );
NAND2_X2 inst_4197 ( .ZN(net_5301), .A1(net_5059), .A2(net_5058) );
CLKBUF_X2 inst_15784 ( .A(net_15631), .Z(net_15632) );
CLKBUF_X2 inst_16151 ( .A(net_15998), .Z(net_15999) );
CLKBUF_X2 inst_15914 ( .A(net_15761), .Z(net_15762) );
CLKBUF_X2 inst_15354 ( .A(net_10840), .Z(net_15202) );
DFFR_X1 inst_7400 ( .D(net_5723), .CK(net_14056), .RN(x6501), .Q(x352) );
CLKBUF_X2 inst_13745 ( .A(net_13592), .Z(net_13593) );
CLKBUF_X2 inst_17176 ( .A(net_17023), .Z(net_17024) );
NAND2_X2 inst_4524 ( .A1(net_3573), .ZN(net_3565), .A2(net_3563) );
NAND2_X2 inst_4871 ( .A1(net_2551), .ZN(net_1158), .A2(net_818) );
CLKBUF_X2 inst_16030 ( .A(net_15877), .Z(net_15878) );
INV_X4 inst_5520 ( .A(net_917), .ZN(net_673) );
NAND2_X2 inst_4257 ( .A1(net_6910), .A2(net_5247), .ZN(net_5203) );
NAND2_X2 inst_4586 ( .A2(net_2947), .ZN(net_2907), .A1(net_2906) );
CLKBUF_X2 inst_18342 ( .A(net_12080), .Z(net_18190) );
CLKBUF_X2 inst_13722 ( .A(net_9796), .Z(net_13570) );
SDFF_X2 inst_1317 ( .Q(net_8087), .D(net_8087), .SE(net_2707), .SI(net_2573), .CK(net_18086) );
DFF_X1 inst_6820 ( .QN(net_8234), .D(net_4447), .CK(net_17204) );
CLKBUF_X2 inst_9623 ( .A(net_9068), .Z(net_9471) );
CLKBUF_X2 inst_12603 ( .A(net_12450), .Z(net_12451) );
SDFF_X2 inst_624 ( .SI(net_8536), .Q(net_8536), .SE(net_3979), .D(net_3967), .CK(net_10159) );
INV_X2 inst_6284 ( .ZN(net_4217), .A(net_3930) );
CLKBUF_X2 inst_17767 ( .A(net_17614), .Z(net_17615) );
INV_X4 inst_5728 ( .A(net_7245), .ZN(net_1955) );
INV_X2 inst_6404 ( .ZN(net_1111), .A(net_1110) );
INV_X2 inst_6419 ( .ZN(net_779), .A(net_778) );
CLKBUF_X2 inst_9886 ( .A(net_9733), .Z(net_9734) );
CLKBUF_X2 inst_18327 ( .A(net_18174), .Z(net_18175) );
CLKBUF_X2 inst_11247 ( .A(net_11094), .Z(net_11095) );
CLKBUF_X2 inst_9375 ( .A(net_9222), .Z(net_9223) );
NAND4_X4 inst_3624 ( .A4(net_3170), .ZN(net_2961), .A2(net_2663), .A1(net_2662), .A3(net_480) );
CLKBUF_X2 inst_17048 ( .A(net_16895), .Z(net_16896) );
CLKBUF_X2 inst_13207 ( .A(net_13054), .Z(net_13055) );
CLKBUF_X2 inst_14598 ( .A(net_14445), .Z(net_14446) );
CLKBUF_X2 inst_11440 ( .A(net_11287), .Z(net_11288) );
CLKBUF_X2 inst_12389 ( .A(net_12236), .Z(net_12237) );
CLKBUF_X2 inst_16495 ( .A(net_10064), .Z(net_16343) );
CLKBUF_X2 inst_13262 ( .A(net_13109), .Z(net_13110) );
CLKBUF_X2 inst_14805 ( .A(net_14652), .Z(net_14653) );
NAND2_X2 inst_4532 ( .A1(net_3381), .ZN(net_3380), .A2(net_3373) );
INV_X2 inst_6277 ( .ZN(net_4271), .A(net_4229) );
CLKBUF_X2 inst_12962 ( .A(net_12809), .Z(net_12810) );
INV_X4 inst_5600 ( .A(net_7362), .ZN(net_1936) );
NOR2_X2 inst_3508 ( .A2(net_2400), .A1(net_2389), .ZN(net_2114) );
INV_X4 inst_5132 ( .ZN(net_5588), .A(net_4357) );
INV_X2 inst_6327 ( .ZN(net_3214), .A(net_3184) );
CLKBUF_X2 inst_14955 ( .A(net_14802), .Z(net_14803) );
CLKBUF_X2 inst_18519 ( .A(net_12034), .Z(net_18367) );
SDFF_X2 inst_1133 ( .D(net_7313), .SI(net_6555), .Q(net_6555), .SE(net_3070), .CK(net_11997) );
NAND2_X2 inst_4580 ( .A2(net_4362), .ZN(net_2956), .A1(net_2955) );
CLKBUF_X2 inst_9990 ( .A(net_9837), .Z(net_9838) );
SDFFR_X2 inst_2103 ( .SE(net_5942), .SI(net_5941), .Q(net_387), .D(net_387), .CK(net_14724), .RN(x6501) );
CLKBUF_X2 inst_16577 ( .A(net_16424), .Z(net_16425) );
AOI221_X4 inst_8710 ( .C1(net_7935), .B1(net_7833), .C2(net_6103), .ZN(net_6043), .B2(net_4398), .A(net_4291) );
CLKBUF_X2 inst_14040 ( .A(net_13887), .Z(net_13888) );
CLKBUF_X2 inst_16234 ( .A(net_16081), .Z(net_16082) );
XNOR2_X2 inst_339 ( .A(net_7388), .ZN(net_783), .B(net_197) );
NAND2_X2 inst_4750 ( .ZN(net_2721), .A1(net_1778), .A2(net_1586) );
CLKBUF_X2 inst_17551 ( .A(net_15319), .Z(net_17399) );
CLKBUF_X2 inst_13995 ( .A(net_13842), .Z(net_13843) );
SDFF_X2 inst_351 ( .SI(net_8463), .Q(net_8463), .SE(net_3983), .D(net_3958), .CK(net_10947) );
CLKBUF_X2 inst_17379 ( .A(net_17226), .Z(net_17227) );
INV_X2 inst_6615 ( .A(net_6209), .ZN(net_6208) );
CLKBUF_X2 inst_10257 ( .A(net_10006), .Z(net_10105) );
CLKBUF_X2 inst_9557 ( .A(net_9404), .Z(net_9405) );
AOI22_X2 inst_7852 ( .A2(net_5595), .ZN(net_4655), .B2(net_4388), .B1(net_2592), .A1(net_322) );
CLKBUF_X2 inst_12507 ( .A(net_12354), .Z(net_12355) );
SDFF_X2 inst_1560 ( .Q(net_7899), .D(net_7899), .SI(net_2711), .SE(net_2543), .CK(net_17001) );
CLKBUF_X2 inst_11463 ( .A(net_11310), .Z(net_11311) );
CLKBUF_X2 inst_12622 ( .A(net_10104), .Z(net_12470) );
CLKBUF_X2 inst_10868 ( .A(net_10715), .Z(net_10716) );
CLKBUF_X2 inst_10994 ( .A(net_9449), .Z(net_10842) );
CLKBUF_X2 inst_13915 ( .A(net_9781), .Z(net_13763) );
CLKBUF_X2 inst_10203 ( .A(net_9764), .Z(net_10051) );
DFFR_X2 inst_7035 ( .QN(net_7492), .D(net_5040), .CK(net_16588), .RN(x6501) );
CLKBUF_X2 inst_9224 ( .A(net_9071), .Z(net_9072) );
CLKBUF_X2 inst_15205 ( .A(net_15052), .Z(net_15053) );
CLKBUF_X2 inst_11164 ( .A(net_11011), .Z(net_11012) );
CLKBUF_X2 inst_10161 ( .A(net_9299), .Z(net_10009) );
SDFF_X2 inst_847 ( .SI(net_8632), .Q(net_8632), .D(net_3980), .SE(net_3885), .CK(net_13323) );
SDFFR_X1 inst_2720 ( .SI(net_9030), .Q(net_9030), .D(net_7459), .SE(net_3208), .CK(net_10676), .RN(x6501) );
INV_X2 inst_6577 ( .ZN(net_798), .A(net_218) );
SDFF_X2 inst_1716 ( .Q(net_7984), .D(net_7984), .SI(net_2702), .SE(net_2542), .CK(net_15242) );
SDFF_X2 inst_1942 ( .SI(net_8076), .Q(net_8076), .D(net_2656), .SE(net_2508), .CK(net_13999) );
CLKBUF_X2 inst_10857 ( .A(net_10365), .Z(net_10705) );
CLKBUF_X2 inst_18271 ( .A(net_18118), .Z(net_18119) );
CLKBUF_X2 inst_9788 ( .A(net_9626), .Z(net_9636) );
INV_X4 inst_5950 ( .ZN(net_2737), .A(net_275) );
CLKBUF_X2 inst_13573 ( .A(net_13420), .Z(net_13421) );
AND2_X4 inst_9136 ( .ZN(net_1397), .A2(net_799), .A1(net_173) );
SDFFR_X1 inst_2648 ( .D(net_6771), .SE(net_4506), .CK(net_9241), .RN(x6501), .SI(x1745), .Q(x1745) );
DFFR_X2 inst_7055 ( .QN(net_7500), .D(net_4778), .CK(net_16674), .RN(x6501) );
CLKBUF_X2 inst_15470 ( .A(net_12139), .Z(net_15318) );
AOI22_X2 inst_7919 ( .A1(net_8995), .A2(net_5456), .B2(net_5260), .ZN(net_4463), .B1(net_3334) );
AOI22_X2 inst_8372 ( .B1(net_8559), .A1(net_8448), .A2(net_6263), .B2(net_6262), .ZN(net_3676) );
SDFF_X2 inst_1146 ( .SI(net_7326), .Q(net_6601), .D(net_6601), .SE(net_3069), .CK(net_11280) );
CLKBUF_X2 inst_18503 ( .A(net_18350), .Z(net_18351) );
CLKBUF_X2 inst_12947 ( .A(net_12794), .Z(net_12795) );
NAND4_X2 inst_3708 ( .A4(net_6222), .A1(net_6221), .ZN(net_4429), .A2(net_3713), .A3(net_3712) );
CLKBUF_X2 inst_18570 ( .A(net_18417), .Z(net_18418) );
NAND2_X4 inst_4023 ( .A1(net_6063), .ZN(net_5982), .A2(net_2247) );
NAND4_X2 inst_3673 ( .A4(net_6052), .A1(net_6051), .ZN(net_4592), .A2(net_4054), .A3(net_4053) );
OAI21_X2 inst_3105 ( .ZN(net_2503), .B2(net_2502), .A(net_2304), .B1(net_2243) );
INV_X4 inst_5162 ( .A(net_3250), .ZN(net_3248) );
CLKBUF_X2 inst_18422 ( .A(net_18269), .Z(net_18270) );
NAND2_X2 inst_4519 ( .ZN(net_3577), .A2(net_3574), .A1(net_3568) );
INV_X4 inst_5349 ( .ZN(net_1724), .A(net_1371) );
INV_X2 inst_6210 ( .ZN(net_5500), .A(net_5389) );
CLKBUF_X2 inst_9899 ( .A(net_9746), .Z(net_9747) );
NOR2_X2 inst_3539 ( .ZN(net_2768), .A1(net_1500), .A2(net_1374) );
SDFFR_X2 inst_2457 ( .QN(net_7412), .SE(net_3354), .SI(net_1457), .CK(net_10093), .D(x13994), .RN(x6501) );
CLKBUF_X2 inst_16442 ( .A(net_12437), .Z(net_16290) );
AOI22_X2 inst_8307 ( .B1(net_8770), .A1(net_8400), .A2(net_3867), .B2(net_3866), .ZN(net_3738) );
CLKBUF_X2 inst_10188 ( .A(net_10035), .Z(net_10036) );
XNOR2_X2 inst_274 ( .A(net_7577), .B(net_3009), .ZN(net_1035) );
CLKBUF_X2 inst_15076 ( .A(net_14810), .Z(net_14924) );
CLKBUF_X2 inst_14543 ( .A(net_14390), .Z(net_14391) );
DFFR_X2 inst_7329 ( .D(net_6825), .QN(net_6822), .CK(net_17929), .RN(x6501) );
OR2_X4 inst_2817 ( .ZN(net_4508), .A2(net_4472), .A1(net_4389) );
CLKBUF_X2 inst_13135 ( .A(net_12982), .Z(net_12983) );
CLKBUF_X2 inst_13436 ( .A(net_13110), .Z(net_13284) );
OAI211_X2 inst_3207 ( .B(net_8903), .ZN(net_2427), .C1(net_2093), .C2(net_2003), .A(net_1059) );
OAI21_X2 inst_3143 ( .B2(net_2060), .ZN(net_2052), .A(net_1985), .B1(net_1681) );
DFFR_X2 inst_7112 ( .QN(net_7607), .D(net_3067), .CK(net_9814), .RN(x6501) );
CLKBUF_X2 inst_11387 ( .A(net_11234), .Z(net_11235) );
SDFFR_X1 inst_2696 ( .SI(net_7529), .SE(net_5043), .CK(net_11947), .RN(x6501), .Q(x4192), .D(x4192) );
CLKBUF_X2 inst_14063 ( .A(net_10308), .Z(net_13911) );
DFFR_X2 inst_7136 ( .QN(net_9050), .D(net_3004), .CK(net_13527), .RN(x6501) );
OR2_X2 inst_2880 ( .ZN(net_2583), .A1(net_2582), .A2(net_2386) );
SDFF_X2 inst_1771 ( .SI(net_6996), .Q(net_6996), .SE(net_6283), .D(net_2544), .CK(net_15888) );
CLKBUF_X2 inst_14402 ( .A(net_14249), .Z(net_14250) );
SDFFR_X1 inst_2660 ( .D(net_6782), .SE(net_4506), .CK(net_11409), .RN(x6501), .SI(x1383), .Q(x1383) );
AOI22_X2 inst_7859 ( .B2(net_5260), .ZN(net_4648), .A2(net_4647), .B1(net_2935), .A1(net_302) );
CLKBUF_X2 inst_13729 ( .A(net_13576), .Z(net_13577) );
SDFFR_X2 inst_2389 ( .SE(net_2260), .Q(net_366), .D(net_366), .CK(net_11450), .RN(x6501), .SI(x1778) );
CLKBUF_X2 inst_17967 ( .A(net_17814), .Z(net_17815) );
INV_X4 inst_5912 ( .A(net_7590), .ZN(net_714) );
CLKBUF_X2 inst_10802 ( .A(net_10649), .Z(net_10650) );
CLKBUF_X2 inst_16906 ( .A(net_16753), .Z(net_16754) );
INV_X2 inst_6199 ( .ZN(net_5511), .A(net_5433) );
CLKBUF_X2 inst_16406 ( .A(net_16253), .Z(net_16254) );
MUX2_X2 inst_4946 ( .B(net_6166), .S(net_3354), .Z(net_2509), .A(x13271) );
SDFFR_X2 inst_2148 ( .QN(net_8262), .SE(net_2996), .D(net_2993), .SI(net_2029), .CK(net_18459), .RN(x6501) );
INV_X4 inst_5784 ( .A(net_7591), .ZN(net_547) );
CLKBUF_X2 inst_17947 ( .A(net_17794), .Z(net_17795) );
CLKBUF_X2 inst_13488 ( .A(net_13134), .Z(net_13336) );
OR2_X2 inst_2900 ( .ZN(net_1304), .A2(x13969), .A1(x13950) );
NOR4_X2 inst_3247 ( .ZN(net_1555), .A3(net_1048), .A4(net_1046), .A2(net_1035), .A1(net_982) );
CLKBUF_X2 inst_13544 ( .A(net_12614), .Z(net_13392) );
SDFF_X2 inst_379 ( .SI(net_8402), .Q(net_8402), .SE(net_3969), .D(net_3951), .CK(net_13440) );
SDFF_X2 inst_926 ( .SI(net_8735), .Q(net_8735), .SE(net_6195), .D(net_3951), .CK(net_11121) );
CLKBUF_X2 inst_12348 ( .A(net_12041), .Z(net_12196) );
CLKBUF_X2 inst_10997 ( .A(net_10688), .Z(net_10845) );
NAND2_X2 inst_4153 ( .ZN(net_5363), .A2(net_5208), .A1(net_5102) );
CLKBUF_X2 inst_13586 ( .A(net_13433), .Z(net_13434) );
AOI222_X1 inst_8684 ( .B1(net_6483), .A2(net_3296), .B2(net_3295), .C2(net_3294), .ZN(net_3288), .A1(net_3282), .C1(net_1542) );
CLKBUF_X2 inst_10624 ( .A(net_9854), .Z(net_10472) );
CLKBUF_X2 inst_15741 ( .A(net_15588), .Z(net_15589) );
CLKBUF_X2 inst_16884 ( .A(net_14436), .Z(net_16732) );
NAND4_X2 inst_3646 ( .ZN(net_4915), .A3(net_4654), .A2(net_4525), .A4(net_4524), .A1(net_4461) );
SDFF_X2 inst_891 ( .Q(net_8575), .D(net_8575), .SI(net_3974), .SE(net_3878), .CK(net_12237) );
CLKBUF_X2 inst_9479 ( .A(net_9140), .Z(net_9327) );
INV_X4 inst_5682 ( .ZN(net_2692), .A(net_276) );
XNOR2_X2 inst_288 ( .B(net_7377), .ZN(net_1006), .A(net_481) );
CLKBUF_X2 inst_14414 ( .A(net_14261), .Z(net_14262) );
CLKBUF_X2 inst_11729 ( .A(net_10155), .Z(net_11577) );
DFFR_X2 inst_7263 ( .QN(net_7402), .D(net_1971), .CK(net_17858), .RN(x6501) );
SDFF_X2 inst_1298 ( .Q(net_7817), .D(net_7817), .SE(net_2730), .SI(net_2706), .CK(net_18089) );
CLKBUF_X2 inst_15059 ( .A(net_14906), .Z(net_14907) );
CLKBUF_X2 inst_14636 ( .A(net_14483), .Z(net_14484) );
AND2_X4 inst_9147 ( .ZN(net_1298), .A2(net_225), .A1(net_181) );
CLKBUF_X2 inst_14856 ( .A(net_12825), .Z(net_14704) );
CLKBUF_X2 inst_12032 ( .A(net_9574), .Z(net_11880) );
AOI22_X2 inst_8241 ( .B1(net_8557), .A1(net_8446), .A2(net_6263), .B2(net_6262), .ZN(net_3796) );
INV_X2 inst_6499 ( .A(net_7434), .ZN(net_544) );
CLKBUF_X2 inst_18484 ( .A(net_13763), .Z(net_18332) );
SDFF_X2 inst_372 ( .SI(net_8538), .Q(net_8538), .SE(net_3979), .D(net_3974), .CK(net_10042) );
DFFR_X1 inst_7388 ( .D(net_5858), .CK(net_14063), .RN(x6501), .Q(x420) );
AOI22_X2 inst_8031 ( .A1(net_7965), .B1(net_7795), .A2(net_6092), .B2(net_6091), .ZN(net_4107) );
CLKBUF_X2 inst_15142 ( .A(net_14989), .Z(net_14990) );
CLKBUF_X2 inst_14623 ( .A(net_14470), .Z(net_14471) );
CLKBUF_X2 inst_9218 ( .A(net_9065), .Z(net_9066) );
AOI22_X2 inst_8512 ( .B1(net_6550), .A1(net_6517), .A2(net_6137), .B2(net_6104), .ZN(net_3428) );
INV_X4 inst_5835 ( .A(net_8256), .ZN(net_1206) );
CLKBUF_X2 inst_11128 ( .A(net_10975), .Z(net_10976) );
SDFF_X2 inst_1775 ( .D(net_7302), .SI(net_6999), .Q(net_6999), .SE(net_6283), .CK(net_18597) );
INV_X2 inst_6223 ( .ZN(net_5487), .A(net_5337) );
SDFF_X2 inst_1172 ( .D(net_7333), .SI(net_6509), .Q(net_6509), .SE(net_3071), .CK(net_18615) );
NAND3_X2 inst_3903 ( .ZN(net_5635), .A1(net_5564), .A3(net_5498), .A2(net_5382) );
CLKBUF_X2 inst_17606 ( .A(net_17453), .Z(net_17454) );
DFFR_X1 inst_7467 ( .QN(net_7443), .D(net_4326), .CK(net_12936), .RN(x6501) );
CLKBUF_X2 inst_13454 ( .A(net_13301), .Z(net_13302) );
CLKBUF_X2 inst_17400 ( .A(net_10496), .Z(net_17248) );
SDFF_X2 inst_1239 ( .Q(net_7834), .D(net_7834), .SE(net_2730), .SI(net_2715), .CK(net_14195) );
CLKBUF_X2 inst_18583 ( .A(net_13584), .Z(net_18431) );
AOI21_X2 inst_8991 ( .B1(net_7526), .ZN(net_1502), .B2(net_1501), .A(net_1354) );
CLKBUF_X2 inst_13832 ( .A(net_13679), .Z(net_13680) );
CLKBUF_X2 inst_14068 ( .A(net_13915), .Z(net_13916) );
DFFR_X2 inst_7094 ( .Q(net_6459), .D(net_3346), .CK(net_15115), .RN(x6501) );
CLKBUF_X2 inst_17468 ( .A(net_17315), .Z(net_17316) );
CLKBUF_X2 inst_11319 ( .A(net_11166), .Z(net_11167) );
AOI22_X2 inst_8556 ( .B2(net_4889), .A1(net_4803), .ZN(net_2917), .B1(net_2916), .A2(net_2568) );
CLKBUF_X2 inst_17427 ( .A(net_17274), .Z(net_17275) );
CLKBUF_X2 inst_14445 ( .A(net_14292), .Z(net_14293) );
AOI22_X2 inst_8300 ( .B1(net_8695), .A1(net_8658), .B2(net_6109), .A2(net_3857), .ZN(net_3743) );
CLKBUF_X2 inst_18199 ( .A(net_18046), .Z(net_18047) );
CLKBUF_X2 inst_13235 ( .A(net_13082), .Z(net_13083) );
CLKBUF_X2 inst_10580 ( .A(net_10427), .Z(net_10428) );
AOI21_X2 inst_8907 ( .ZN(net_5795), .A(net_5745), .B2(net_5606), .B1(net_4910) );
INV_X4 inst_5088 ( .ZN(net_5711), .A(net_5687) );
CLKBUF_X2 inst_16938 ( .A(net_16785), .Z(net_16786) );
NAND2_X2 inst_4193 ( .ZN(net_5306), .A1(net_5181), .A2(net_4983) );
CLKBUF_X2 inst_17287 ( .A(net_17134), .Z(net_17135) );
CLKBUF_X2 inst_13316 ( .A(net_9952), .Z(net_13164) );
DFFR_X2 inst_7074 ( .D(net_3925), .QN(net_476), .CK(net_11246), .RN(x6501) );
CLKBUF_X2 inst_14200 ( .A(net_13754), .Z(net_14048) );
CLKBUF_X2 inst_12858 ( .A(net_12705), .Z(net_12706) );
SDFF_X2 inst_686 ( .Q(net_8677), .D(net_8677), .SI(net_3960), .SE(net_3935), .CK(net_11071) );
CLKBUF_X2 inst_9871 ( .A(net_9718), .Z(net_9719) );
CLKBUF_X2 inst_14777 ( .A(net_14624), .Z(net_14625) );
NAND2_X2 inst_4892 ( .A2(net_7379), .ZN(net_700), .A1(net_168) );
NAND4_X2 inst_3643 ( .ZN(net_4918), .A4(net_4649), .A3(net_4565), .A2(net_4520), .A1(net_4499) );
CLKBUF_X2 inst_10635 ( .A(net_10482), .Z(net_10483) );
AND2_X4 inst_9075 ( .ZN(net_3247), .A1(net_3177), .A2(net_3176) );
SDFFR_X2 inst_2119 ( .SI(net_7194), .Q(net_7194), .D(net_6445), .SE(net_4362), .CK(net_13574), .RN(x6501) );
SDFF_X2 inst_1929 ( .SI(net_8056), .Q(net_8056), .D(net_2574), .SE(net_2508), .CK(net_16023) );
NOR2_X2 inst_3391 ( .ZN(net_4834), .A2(net_4473), .A1(net_1432) );
CLKBUF_X2 inst_9422 ( .A(net_9269), .Z(net_9270) );
AOI22_X2 inst_8519 ( .B1(net_6618), .A1(net_6585), .A2(net_6257), .B2(net_6110), .ZN(net_3421) );
AND4_X4 inst_9025 ( .ZN(net_4969), .A4(net_4720), .A1(net_4577), .A2(net_4539), .A3(net_4481) );
CLKBUF_X2 inst_12472 ( .A(net_12319), .Z(net_12320) );
SDFF_X2 inst_1794 ( .D(net_7278), .SI(net_6935), .Q(net_6935), .SE(net_6281), .CK(net_14627) );
CLKBUF_X2 inst_15023 ( .A(net_14870), .Z(net_14871) );
AOI22_X2 inst_8126 ( .B1(net_8151), .A1(net_7709), .B2(net_6101), .A2(net_6095), .ZN(net_6028) );
CLKBUF_X2 inst_16010 ( .A(net_9888), .Z(net_15858) );
OAI21_X2 inst_3047 ( .B2(net_8244), .B1(net_4954), .ZN(net_4772), .A(net_4497) );
INV_X4 inst_5957 ( .ZN(net_518), .A(x494) );
NAND4_X2 inst_3847 ( .ZN(net_2304), .A3(net_1936), .A4(net_1750), .A1(net_1293), .A2(net_1056) );
CLKBUF_X2 inst_18464 ( .A(net_9719), .Z(net_18312) );
CLKBUF_X2 inst_14494 ( .A(net_14341), .Z(net_14342) );
CLKBUF_X2 inst_18192 ( .A(net_18039), .Z(net_18040) );
INV_X4 inst_5756 ( .A(net_6296), .ZN(net_630) );
CLKBUF_X2 inst_11376 ( .A(net_11223), .Z(net_11224) );
CLKBUF_X2 inst_14369 ( .A(net_14216), .Z(net_14217) );
CLKBUF_X2 inst_9748 ( .A(net_9072), .Z(net_9596) );
SDFF_X2 inst_1660 ( .SI(net_7751), .Q(net_7751), .D(net_2720), .SE(net_2560), .CK(net_18361) );
CLKBUF_X2 inst_10113 ( .A(net_9320), .Z(net_9961) );
NAND2_X2 inst_4375 ( .A1(net_7115), .A2(net_5164), .ZN(net_5082) );
CLKBUF_X2 inst_13416 ( .A(net_10565), .Z(net_13264) );
SDFF_X2 inst_517 ( .Q(net_8871), .D(net_8871), .SI(net_3974), .SE(net_3936), .CK(net_12277) );
SDFF_X2 inst_1261 ( .Q(net_8106), .D(net_8106), .SI(net_2715), .SE(net_2707), .CK(net_14297) );
INV_X4 inst_5368 ( .A(net_1962), .ZN(net_1133) );
AOI21_X2 inst_8967 ( .B1(net_7645), .B2(net_6181), .ZN(net_3005), .A(net_2533) );
CLKBUF_X2 inst_10220 ( .A(net_10067), .Z(net_10068) );
INV_X4 inst_6130 ( .A(net_6333), .ZN(net_757) );
INV_X4 inst_5382 ( .ZN(net_2785), .A(net_1363) );
CLKBUF_X2 inst_14661 ( .A(net_14508), .Z(net_14509) );
XNOR2_X2 inst_310 ( .B(net_2150), .ZN(net_961), .A(net_586) );
CLKBUF_X2 inst_18875 ( .A(net_18722), .Z(net_18723) );
CLKBUF_X2 inst_17982 ( .A(net_17829), .Z(net_17830) );
AOI21_X2 inst_8900 ( .B2(net_5871), .ZN(net_5780), .A(net_5762), .B1(x275) );
SDFFR_X1 inst_2688 ( .SI(net_7551), .SE(net_5043), .CK(net_12752), .RN(x6501), .Q(x3904), .D(x3904) );
INV_X32 inst_6172 ( .ZN(net_5016), .A(net_4709) );
INV_X4 inst_5592 ( .A(net_8954), .ZN(net_1271) );
CLKBUF_X2 inst_18091 ( .A(net_17938), .Z(net_17939) );
SDFFR_X2 inst_2351 ( .SE(net_2260), .Q(net_313), .D(net_313), .CK(net_10464), .RN(x6501), .SI(x3418) );
AOI22_X2 inst_8067 ( .B1(net_8140), .A1(net_7902), .A2(net_6098), .B2(net_4190), .ZN(net_4076) );
CLKBUF_X2 inst_12302 ( .A(net_12149), .Z(net_12150) );
INV_X4 inst_5125 ( .ZN(net_5267), .A(net_4395) );
SDFF_X2 inst_1853 ( .D(net_7277), .SI(net_6934), .Q(net_6934), .SE(net_6281), .CK(net_17355) );
DFFR_X1 inst_7576 ( .Q(net_8285), .D(net_8275), .CK(net_12226), .RN(x6501) );
CLKBUF_X2 inst_11101 ( .A(net_10948), .Z(net_10949) );
XNOR2_X2 inst_264 ( .B(net_6831), .A(net_1221), .ZN(net_1120) );
CLKBUF_X2 inst_15834 ( .A(net_15681), .Z(net_15682) );
NAND4_X2 inst_3710 ( .A4(net_6238), .A1(net_6237), .ZN(net_4427), .A2(net_3700), .A3(net_3699) );
SDFF_X2 inst_1260 ( .Q(net_8104), .D(net_8104), .SI(net_2710), .SE(net_2707), .CK(net_14443) );
INV_X2 inst_6490 ( .A(net_6472), .ZN(net_3286) );
CLKBUF_X2 inst_10190 ( .A(net_10037), .Z(net_10038) );
NOR2_X4 inst_3332 ( .ZN(net_6186), .A1(net_6143), .A2(net_3079) );
AOI22_X2 inst_7885 ( .B1(net_8996), .A2(net_5538), .B2(net_5456), .ZN(net_4546), .A1(net_425) );
NAND2_X2 inst_4898 ( .A2(net_7390), .ZN(net_639), .A1(net_179) );
CLKBUF_X2 inst_17126 ( .A(net_16973), .Z(net_16974) );
SDFFR_X1 inst_2717 ( .SI(net_9026), .Q(net_9026), .D(net_7455), .SE(net_3208), .CK(net_12846), .RN(x6501) );
CLKBUF_X2 inst_13836 ( .A(net_13683), .Z(net_13684) );
NAND2_X2 inst_4176 ( .ZN(net_5330), .A1(net_5080), .A2(net_5079) );
XNOR2_X2 inst_129 ( .ZN(net_2825), .A(net_2552), .B(net_818) );
SDFFR_X1 inst_2740 ( .SI(net_9023), .Q(net_9023), .D(net_7452), .SE(net_3208), .CK(net_10095), .RN(x6501) );
SDFF_X2 inst_1754 ( .SI(net_7739), .Q(net_7739), .D(net_2585), .SE(net_2560), .CK(net_15739) );
CLKBUF_X2 inst_16777 ( .A(net_16624), .Z(net_16625) );
DFFR_X2 inst_6974 ( .QN(net_5965), .D(net_5917), .CK(net_9285), .RN(x6501) );
CLKBUF_X2 inst_12955 ( .A(net_12802), .Z(net_12803) );
AOI22_X2 inst_7789 ( .A2(net_6187), .B2(net_5463), .ZN(net_4811), .B1(net_436), .A1(net_199) );
SDFFR_X1 inst_2727 ( .SI(net_9039), .Q(net_9039), .D(net_7468), .SE(net_3208), .CK(net_10657), .RN(x6501) );
AOI22_X2 inst_7974 ( .B1(net_8094), .A1(net_7754), .B2(net_6108), .A2(net_6096), .ZN(net_4156) );
AOI221_X2 inst_8848 ( .B1(net_8866), .C1(net_8311), .B2(net_6252), .ZN(net_6245), .C2(net_4345), .A(net_4262) );
INV_X2 inst_6305 ( .ZN(net_3899), .A(net_3601) );
CLKBUF_X2 inst_18664 ( .A(net_18511), .Z(net_18512) );
SDFF_X2 inst_777 ( .SI(net_8345), .Q(net_8345), .D(net_3962), .SE(net_3880), .CK(net_12424) );
INV_X4 inst_6164 ( .A(net_6272), .ZN(net_6271) );
CLKBUF_X2 inst_14175 ( .A(net_12255), .Z(net_14023) );
INV_X8 inst_5016 ( .ZN(net_5655), .A(net_4386) );
CLKBUF_X2 inst_17872 ( .A(net_17719), .Z(net_17720) );
CLKBUF_X2 inst_17199 ( .A(net_12230), .Z(net_17047) );
CLKBUF_X2 inst_10276 ( .A(net_10123), .Z(net_10124) );
DFFR_X2 inst_7000 ( .QN(net_5960), .D(net_5874), .CK(net_9276), .RN(x6501) );
CLKBUF_X2 inst_15975 ( .A(net_15822), .Z(net_15823) );
CLKBUF_X2 inst_9983 ( .A(net_9643), .Z(net_9831) );
NAND4_X2 inst_3724 ( .ZN(net_4306), .A1(net_4172), .A2(net_4171), .A3(net_4170), .A4(net_4169) );
CLKBUF_X2 inst_14393 ( .A(net_14240), .Z(net_14241) );
CLKBUF_X2 inst_14138 ( .A(net_13985), .Z(net_13986) );
CLKBUF_X2 inst_15943 ( .A(net_15790), .Z(net_15791) );
CLKBUF_X2 inst_16930 ( .A(net_14653), .Z(net_16778) );
CLKBUF_X2 inst_10509 ( .A(net_10356), .Z(net_10357) );
INV_X4 inst_6146 ( .A(net_6806), .ZN(net_6140) );
CLKBUF_X2 inst_13978 ( .A(net_13825), .Z(net_13826) );
CLKBUF_X2 inst_11909 ( .A(net_11756), .Z(net_11757) );
MUX2_X2 inst_4965 ( .A(net_7389), .S(net_2370), .Z(net_2358), .B(net_795) );
CLKBUF_X2 inst_13039 ( .A(net_11283), .Z(net_12887) );
CLKBUF_X2 inst_11158 ( .A(net_11005), .Z(net_11006) );
SDFFR_X2 inst_2354 ( .QN(net_7479), .SE(net_3354), .SI(net_3127), .CK(net_9965), .D(x13341), .RN(x6501) );
CLKBUF_X2 inst_9447 ( .A(net_9294), .Z(net_9295) );
AOI221_X4 inst_8735 ( .B1(net_8818), .C1(net_8337), .C2(net_6265), .B2(net_6253), .ZN(net_4331), .A(net_4237) );
CLKBUF_X2 inst_10729 ( .A(net_10576), .Z(net_10577) );
CLKBUF_X2 inst_13315 ( .A(net_13162), .Z(net_13163) );
CLKBUF_X2 inst_15514 ( .A(net_9519), .Z(net_15362) );
CLKBUF_X2 inst_15872 ( .A(net_15719), .Z(net_15720) );
CLKBUF_X2 inst_14965 ( .A(net_14812), .Z(net_14813) );
CLKBUF_X2 inst_12316 ( .A(net_12163), .Z(net_12164) );
CLKBUF_X2 inst_10883 ( .A(net_10730), .Z(net_10731) );
NAND3_X4 inst_3869 ( .A1(net_6261), .A3(net_6190), .A2(net_4816), .ZN(net_4814) );
NOR2_X2 inst_3488 ( .ZN(net_2220), .A1(net_2093), .A2(net_1889) );
CLKBUF_X2 inst_15801 ( .A(net_15648), .Z(net_15649) );
CLKBUF_X2 inst_12689 ( .A(net_12536), .Z(net_12537) );
NAND2_X2 inst_4563 ( .ZN(net_3887), .A1(net_3251), .A2(net_3178) );
CLKBUF_X2 inst_17813 ( .A(net_17660), .Z(net_17661) );
INV_X4 inst_5504 ( .A(net_976), .ZN(net_694) );
CLKBUF_X2 inst_19134 ( .A(net_18981), .Z(net_18982) );
DFFR_X1 inst_7453 ( .QN(net_8911), .D(net_4740), .CK(net_14850), .RN(x6501) );
SDFF_X2 inst_1519 ( .Q(net_7887), .D(net_7887), .SI(net_2720), .SE(net_2543), .CK(net_15281) );
DFFR_X2 inst_7243 ( .QN(net_5956), .D(net_2055), .CK(net_15055), .RN(x6501) );
CLKBUF_X2 inst_9936 ( .A(net_9783), .Z(net_9784) );
AOI22_X2 inst_8461 ( .B1(net_6719), .A1(net_6686), .B2(net_6202), .A2(net_3520), .ZN(net_3479) );
MUX2_X2 inst_4989 ( .A(net_9031), .Z(net_3944), .B(net_3009), .S(net_622) );
CLKBUF_X2 inst_16617 ( .A(net_9104), .Z(net_16465) );
CLKBUF_X2 inst_18601 ( .A(net_14883), .Z(net_18449) );
NAND2_X2 inst_4324 ( .A1(net_7081), .A2(net_5164), .ZN(net_5133) );
INV_X4 inst_5746 ( .A(net_7497), .ZN(net_3309) );
INV_X4 inst_5597 ( .A(net_7434), .ZN(net_3167) );
CLKBUF_X2 inst_12705 ( .A(net_11738), .Z(net_12553) );
AOI22_X2 inst_8531 ( .B1(net_6591), .A1(net_6558), .A2(net_6257), .B2(net_6110), .ZN(net_3409) );
CLKBUF_X2 inst_12244 ( .A(net_12091), .Z(net_12092) );
SDFF_X2 inst_1491 ( .SI(net_7278), .Q(net_7095), .D(net_7095), .SE(net_6278), .CK(net_14631) );
AOI22_X2 inst_8070 ( .B1(net_8208), .A1(net_7698), .B2(net_6099), .A2(net_4399), .ZN(net_4073) );
CLKBUF_X2 inst_12747 ( .A(net_12594), .Z(net_12595) );
CLKBUF_X2 inst_15446 ( .A(net_15293), .Z(net_15294) );
SDFFR_X1 inst_2676 ( .SI(net_7540), .SE(net_5043), .CK(net_9711), .RN(x6501), .Q(x4059), .D(x4059) );
AOI22_X2 inst_8566 ( .A1(net_2762), .B2(net_2556), .ZN(net_2201), .A2(net_1909), .B1(net_1908) );
XNOR2_X2 inst_154 ( .ZN(net_2017), .B(net_1734), .A(net_1717) );
CLKBUF_X2 inst_9794 ( .A(net_9641), .Z(net_9642) );
INV_X4 inst_6057 ( .A(net_7257), .ZN(net_1947) );
CLKBUF_X2 inst_12325 ( .A(net_12172), .Z(net_12173) );
CLKBUF_X2 inst_10078 ( .A(net_9106), .Z(net_9926) );
CLKBUF_X2 inst_13427 ( .A(net_13274), .Z(net_13275) );
CLKBUF_X2 inst_10368 ( .A(net_10171), .Z(net_10216) );
NAND2_X2 inst_4240 ( .A1(net_7023), .A2(net_5249), .ZN(net_5220) );
CLKBUF_X2 inst_10813 ( .A(net_10660), .Z(net_10661) );
CLKBUF_X2 inst_12570 ( .A(net_12417), .Z(net_12418) );
SDFF_X2 inst_1790 ( .D(net_7288), .SI(net_6985), .Q(net_6985), .SE(net_6283), .CK(net_17685) );
INV_X2 inst_6621 ( .A(net_6272), .ZN(net_6268) );
CLKBUF_X2 inst_10989 ( .A(net_10484), .Z(net_10837) );
INV_X2 inst_6355 ( .ZN(net_2213), .A(net_2212) );
CLKBUF_X2 inst_13982 ( .A(net_13439), .Z(net_13830) );
CLKBUF_X2 inst_18155 ( .A(net_18002), .Z(net_18003) );
XNOR2_X2 inst_243 ( .B(net_7165), .A(net_2031), .ZN(net_1218) );
SDFF_X2 inst_1378 ( .Q(net_8186), .D(net_8186), .SI(net_2708), .SE(net_2561), .CK(net_18286) );
CLKBUF_X2 inst_14156 ( .A(net_14003), .Z(net_14004) );
CLKBUF_X2 inst_14049 ( .A(net_13896), .Z(net_13897) );
CLKBUF_X2 inst_18521 ( .A(net_18368), .Z(net_18369) );
CLKBUF_X2 inst_16894 ( .A(net_15646), .Z(net_16742) );
CLKBUF_X2 inst_15738 ( .A(net_15585), .Z(net_15586) );
AOI22_X2 inst_8189 ( .B1(net_8865), .A1(net_8310), .B2(net_6252), .A2(net_4345), .ZN(net_3844) );
DFFR_X2 inst_7281 ( .QN(net_6388), .D(net_1731), .CK(net_15661), .RN(x6501) );
CLKBUF_X2 inst_16491 ( .A(net_16338), .Z(net_16339) );
HA_X1 inst_6704 ( .CO(net_6176), .S(net_1775), .B(net_1453), .A(x3418) );
CLKBUF_X2 inst_9501 ( .A(net_9155), .Z(net_9349) );
CLKBUF_X2 inst_16709 ( .A(net_11480), .Z(net_16557) );
AOI221_X2 inst_8799 ( .C2(net_6187), .B2(net_5609), .A(net_4898), .ZN(net_4878), .B1(net_371), .C1(net_195) );
NOR4_X2 inst_3229 ( .ZN(net_2110), .A4(net_1832), .A3(net_1560), .A1(net_983), .A2(net_786) );
NAND2_X2 inst_4135 ( .ZN(net_5387), .A1(net_5122), .A2(net_5121) );
CLKBUF_X2 inst_14459 ( .A(net_14306), .Z(net_14307) );
SDFF_X2 inst_1369 ( .SI(net_7867), .Q(net_7867), .D(net_2639), .SE(net_2558), .CK(net_14023) );
NAND3_X2 inst_3988 ( .ZN(net_1682), .A1(net_1483), .A2(net_989), .A3(net_988) );
INV_X2 inst_6548 ( .A(net_6808), .ZN(net_4619) );
CLKBUF_X2 inst_18548 ( .A(net_18395), .Z(net_18396) );
CLKBUF_X2 inst_15172 ( .A(net_15019), .Z(net_15020) );
CLKBUF_X2 inst_15280 ( .A(net_15127), .Z(net_15128) );
SDFFR_X2 inst_2561 ( .QN(net_6357), .SE(net_2147), .SI(net_1807), .D(net_765), .CK(net_14747), .RN(x6501) );
AOI22_X2 inst_7767 ( .B1(net_6994), .A1(net_6954), .A2(net_5443), .B2(net_5442), .ZN(net_5338) );
AOI22_X2 inst_8495 ( .B1(net_6613), .A1(net_6580), .A2(net_6257), .B2(net_6110), .ZN(net_3445) );
AOI21_X2 inst_8974 ( .A(net_8947), .B2(net_6219), .ZN(net_2482), .B1(net_2264) );
AOI22_X2 inst_8163 ( .B1(net_8704), .A1(net_8482), .ZN(net_6073), .B2(net_4350), .A2(net_4349) );
CLKBUF_X2 inst_13669 ( .A(net_13296), .Z(net_13517) );
CLKBUF_X2 inst_13257 ( .A(net_13104), .Z(net_13105) );
CLKBUF_X2 inst_9583 ( .A(net_9430), .Z(net_9431) );
NAND2_X2 inst_4226 ( .A1(net_7017), .A2(net_5249), .ZN(net_5234) );
CLKBUF_X2 inst_16011 ( .A(net_15858), .Z(net_15859) );
CLKBUF_X2 inst_15847 ( .A(net_15694), .Z(net_15695) );
CLKBUF_X2 inst_9222 ( .A(net_9068), .Z(net_9070) );
CLKBUF_X2 inst_12843 ( .A(net_12690), .Z(net_12691) );
INV_X4 inst_5795 ( .A(net_7612), .ZN(net_2549) );
CLKBUF_X2 inst_12112 ( .A(net_11959), .Z(net_11960) );
SDFFR_X2 inst_2238 ( .Q(net_7458), .D(net_7458), .SE(net_2863), .CK(net_10621), .SI(x13520), .RN(x6501) );
INV_X4 inst_5207 ( .A(net_3354), .ZN(net_3352) );
NAND2_X2 inst_4543 ( .ZN(net_3355), .A1(net_3354), .A2(net_3351) );
INV_X4 inst_5072 ( .ZN(net_5856), .A(net_5810) );
CLKBUF_X2 inst_14347 ( .A(net_14194), .Z(net_14195) );
OAI21_X2 inst_3151 ( .B2(net_1984), .ZN(net_1983), .A(net_1977), .B1(net_761) );
CLKBUF_X2 inst_15312 ( .A(net_15151), .Z(net_15160) );
CLKBUF_X2 inst_13073 ( .A(net_12920), .Z(net_12921) );
CLKBUF_X2 inst_10764 ( .A(net_10611), .Z(net_10612) );
NAND2_X2 inst_4436 ( .A1(net_6873), .A2(net_5016), .ZN(net_4991) );
AOI22_X2 inst_8180 ( .A1(net_8604), .B1(net_8419), .A2(net_3864), .B2(net_3863), .ZN(net_3852) );
CLKBUF_X2 inst_16307 ( .A(net_16154), .Z(net_16155) );
CLKBUF_X2 inst_13042 ( .A(net_12889), .Z(net_12890) );
CLKBUF_X2 inst_14732 ( .A(net_14171), .Z(net_14580) );
INV_X4 inst_5801 ( .A(net_7597), .ZN(net_543) );
CLKBUF_X2 inst_9363 ( .A(net_9210), .Z(net_9211) );
HA_X1 inst_6674 ( .S(net_3169), .CO(net_3168), .A(net_3167), .B(net_3089) );
SDFFR_X2 inst_2259 ( .SE(net_2801), .D(net_2796), .SI(net_200), .Q(net_200), .CK(net_14985), .RN(x6501) );
CLKBUF_X2 inst_12935 ( .A(net_10177), .Z(net_12783) );
INV_X2 inst_6196 ( .ZN(net_5514), .A(net_5447) );
CLKBUF_X2 inst_14314 ( .A(net_14161), .Z(net_14162) );
INV_X2 inst_6462 ( .A(net_6412), .ZN(net_580) );
CLKBUF_X2 inst_14101 ( .A(net_12010), .Z(net_13949) );
CLKBUF_X2 inst_12824 ( .A(net_12671), .Z(net_12672) );
CLKBUF_X2 inst_11915 ( .A(net_10384), .Z(net_11763) );
CLKBUF_X2 inst_18232 ( .A(net_18079), .Z(net_18080) );
CLKBUF_X2 inst_12280 ( .A(net_12127), .Z(net_12128) );
CLKBUF_X2 inst_11072 ( .A(net_10919), .Z(net_10920) );
INV_X2 inst_6428 ( .ZN(net_728), .A(net_727) );
CLKBUF_X2 inst_14221 ( .A(net_14068), .Z(net_14069) );
DFFR_X2 inst_7312 ( .D(net_294), .QN(net_153), .CK(net_11136), .RN(x6501) );
CLKBUF_X2 inst_19049 ( .A(net_18896), .Z(net_18897) );
CLKBUF_X2 inst_17731 ( .A(net_17578), .Z(net_17579) );
CLKBUF_X2 inst_17409 ( .A(net_15059), .Z(net_17257) );
CLKBUF_X2 inst_10749 ( .A(net_10596), .Z(net_10597) );
CLKBUF_X2 inst_18479 ( .A(net_17715), .Z(net_18327) );
CLKBUF_X2 inst_12737 ( .A(net_12192), .Z(net_12585) );
CLKBUF_X2 inst_17499 ( .A(net_17346), .Z(net_17347) );
SDFF_X2 inst_524 ( .Q(net_8880), .D(net_8880), .SI(net_3953), .SE(net_3936), .CK(net_10277) );
CLKBUF_X2 inst_15568 ( .A(net_11200), .Z(net_15416) );
CLKBUF_X2 inst_13027 ( .A(net_11592), .Z(net_12875) );
XOR2_X1 inst_104 ( .Z(net_1024), .A(net_1023), .B(net_187) );
CLKBUF_X2 inst_14986 ( .A(net_11392), .Z(net_14834) );
SDFFR_X2 inst_2331 ( .SE(net_2260), .Q(net_338), .D(net_338), .CK(net_11461), .RN(x6501), .SI(x2261) );
INV_X4 inst_6096 ( .A(net_7366), .ZN(net_1778) );
CLKBUF_X2 inst_9752 ( .A(net_9560), .Z(net_9600) );
SDFFR_X2 inst_2377 ( .SE(net_2260), .Q(net_326), .D(net_326), .CK(net_10428), .RN(x6501), .SI(x2856) );
SDFFR_X2 inst_2522 ( .D(net_7371), .SE(net_2387), .SI(net_286), .Q(net_286), .CK(net_16395), .RN(x6501) );
CLKBUF_X2 inst_13793 ( .A(net_10013), .Z(net_13641) );
CLKBUF_X2 inst_11910 ( .A(net_10201), .Z(net_11758) );
CLKBUF_X2 inst_10673 ( .A(net_10520), .Z(net_10521) );
CLKBUF_X2 inst_18530 ( .A(net_18377), .Z(net_18378) );
AOI22_X2 inst_7967 ( .A1(net_7957), .B1(net_7787), .A2(net_6092), .B2(net_6091), .ZN(net_4162) );
INV_X4 inst_5216 ( .ZN(net_2475), .A(net_2323) );
INV_X4 inst_5257 ( .ZN(net_2060), .A(net_1871) );
AOI22_X2 inst_8011 ( .B1(net_8064), .A1(net_7860), .B2(net_6107), .A2(net_4400), .ZN(net_4124) );
CLKBUF_X2 inst_11226 ( .A(net_11073), .Z(net_11074) );
SDFF_X2 inst_708 ( .SI(net_8621), .Q(net_8621), .SE(net_3984), .D(net_3953), .CK(net_10243) );
SDFF_X2 inst_1346 ( .Q(net_8208), .D(net_8208), .SI(net_2715), .SE(net_2561), .CK(net_14186) );
NOR2_X2 inst_3523 ( .A1(net_1910), .ZN(net_1899), .A2(net_1730) );
INV_X4 inst_5811 ( .A(net_6334), .ZN(net_2255) );
NOR2_X2 inst_3510 ( .A1(net_6324), .ZN(net_1838), .A2(net_1837) );
INV_X4 inst_5108 ( .ZN(net_4952), .A(net_4899) );
DFF_X1 inst_6723 ( .Q(net_6769), .D(net_5646), .CK(net_9264) );
SDFF_X2 inst_1071 ( .D(net_7321), .SI(net_6530), .Q(net_6530), .SE(net_3086), .CK(net_12097) );
NAND2_X2 inst_4277 ( .A1(net_6883), .A2(net_5247), .ZN(net_5183) );
INV_X2 inst_6421 ( .ZN(net_766), .A(net_765) );
INV_X4 inst_5291 ( .ZN(net_2077), .A(net_1868) );
CLKBUF_X2 inst_17476 ( .A(net_17323), .Z(net_17324) );
CLKBUF_X2 inst_11352 ( .A(net_9714), .Z(net_11200) );
CLKBUF_X2 inst_17783 ( .A(net_17630), .Z(net_17631) );
CLKBUF_X2 inst_13211 ( .A(net_11074), .Z(net_13059) );
SDFF_X2 inst_1994 ( .SI(net_7938), .Q(net_7938), .D(net_2704), .SE(net_2461), .CK(net_16968) );
CLKBUF_X2 inst_13132 ( .A(net_10937), .Z(net_12980) );
CLKBUF_X2 inst_15952 ( .A(net_15799), .Z(net_15800) );
AND2_X2 inst_9192 ( .A2(net_5691), .ZN(net_1638), .A1(net_1637) );
INV_X4 inst_5298 ( .ZN(net_1773), .A(net_1597) );
CLKBUF_X2 inst_14436 ( .A(net_14283), .Z(net_14284) );
CLKBUF_X2 inst_10108 ( .A(net_9713), .Z(net_9956) );
CLKBUF_X2 inst_15179 ( .A(net_15026), .Z(net_15027) );
CLKBUF_X2 inst_14935 ( .A(net_14782), .Z(net_14783) );
CLKBUF_X2 inst_14744 ( .A(net_14591), .Z(net_14592) );
CLKBUF_X2 inst_13191 ( .A(net_13038), .Z(net_13039) );
AOI21_X2 inst_8940 ( .A(net_5746), .ZN(net_5700), .B2(net_5518), .B1(net_4535) );
SDFFR_X2 inst_2162 ( .QN(net_7580), .D(net_3974), .SE(net_3144), .SI(net_3139), .CK(net_10873), .RN(x6501) );
SDFF_X2 inst_392 ( .Q(net_8826), .D(net_8826), .SE(net_3964), .SI(net_3962), .CK(net_10204) );
XNOR2_X2 inst_120 ( .ZN(net_2984), .A(net_2833), .B(net_1055) );
CLKBUF_X2 inst_14533 ( .A(net_14380), .Z(net_14381) );
AOI22_X2 inst_7747 ( .B1(net_6976), .A1(net_6936), .A2(net_5443), .B2(net_5442), .ZN(net_5418) );
CLKBUF_X2 inst_10917 ( .A(net_9628), .Z(net_10765) );
CLKBUF_X2 inst_17575 ( .A(net_17422), .Z(net_17423) );
SDFF_X2 inst_1514 ( .SI(net_7846), .Q(net_7846), .D(net_2708), .SE(net_2558), .CK(net_18276) );
AOI22_X2 inst_8361 ( .B1(net_8851), .A1(net_8370), .A2(net_6265), .B2(net_6253), .ZN(net_3687) );
SDFF_X2 inst_567 ( .Q(net_8831), .D(net_8831), .SE(net_3964), .SI(net_3944), .CK(net_10842) );
OAI211_X2 inst_3200 ( .ZN(net_2846), .B(net_2329), .A(net_2092), .C1(net_1910), .C2(net_1659) );
AND2_X4 inst_9134 ( .ZN(net_1387), .A2(net_804), .A1(net_172) );
SDFF_X2 inst_1601 ( .Q(net_8136), .D(net_8136), .SI(net_2717), .SE(net_2541), .CK(net_14167) );
NOR2_X2 inst_3526 ( .ZN(net_2070), .A2(net_1701), .A1(net_716) );
AOI211_X2 inst_9010 ( .ZN(net_5532), .C1(net_4926), .A(net_4925), .C2(net_4686), .B(net_3037) );
CLKBUF_X2 inst_18501 ( .A(net_18348), .Z(net_18349) );
CLKBUF_X2 inst_12147 ( .A(net_11994), .Z(net_11995) );
CLKBUF_X2 inst_10910 ( .A(net_10757), .Z(net_10758) );
DFFS_X1 inst_6916 ( .QN(net_6798), .D(net_4682), .CK(net_11809), .SN(x6501) );
CLKBUF_X2 inst_13999 ( .A(net_13846), .Z(net_13847) );
CLKBUF_X2 inst_9876 ( .A(net_9420), .Z(net_9724) );
CLKBUF_X2 inst_18365 ( .A(net_18212), .Z(net_18213) );
NAND2_X2 inst_4123 ( .ZN(net_5403), .A1(net_5134), .A2(net_5133) );
SDFF_X2 inst_1751 ( .SI(net_7768), .Q(net_7768), .D(net_2704), .SE(net_2560), .CK(net_14395) );
DFFS_X1 inst_6919 ( .QN(net_8889), .D(net_3588), .CK(net_11208), .SN(x6501) );
AOI22_X2 inst_7766 ( .B1(net_6993), .A1(net_6953), .A2(net_5443), .B2(net_5442), .ZN(net_5342) );
CLKBUF_X2 inst_14490 ( .A(net_12186), .Z(net_14338) );
AOI22_X2 inst_8140 ( .B1(net_8153), .A1(net_7711), .B2(net_6101), .A2(net_6095), .ZN(net_6032) );
CLKBUF_X2 inst_18388 ( .A(net_18235), .Z(net_18236) );
CLKBUF_X2 inst_17462 ( .A(net_17309), .Z(net_17310) );
SDFFR_X2 inst_2235 ( .QN(net_9055), .SE(net_2963), .SI(net_2827), .D(net_2119), .CK(net_13448), .RN(x6501) );
SDFF_X2 inst_779 ( .SI(net_8347), .Q(net_8347), .D(net_3966), .SE(net_3880), .CK(net_9990) );
CLKBUF_X2 inst_11465 ( .A(net_11312), .Z(net_11313) );
CLKBUF_X2 inst_16563 ( .A(net_16410), .Z(net_16411) );
CLKBUF_X2 inst_18567 ( .A(net_18414), .Z(net_18415) );
CLKBUF_X2 inst_10503 ( .A(net_10350), .Z(net_10351) );
NAND2_X2 inst_4131 ( .ZN(net_5392), .A1(net_5125), .A2(net_5124) );
CLKBUF_X2 inst_17502 ( .A(net_17349), .Z(net_17350) );
CLKBUF_X2 inst_9805 ( .A(net_9652), .Z(net_9653) );
CLKBUF_X2 inst_13591 ( .A(net_13438), .Z(net_13439) );
CLKBUF_X2 inst_18860 ( .A(net_18707), .Z(net_18708) );
CLKBUF_X2 inst_16184 ( .A(net_16031), .Z(net_16032) );
NAND2_X2 inst_4228 ( .A1(net_7018), .A2(net_5249), .ZN(net_5232) );
CLKBUF_X2 inst_15838 ( .A(net_9419), .Z(net_15686) );
CLKBUF_X2 inst_16647 ( .A(net_14114), .Z(net_16495) );
CLKBUF_X2 inst_10808 ( .A(net_9491), .Z(net_10656) );
CLKBUF_X2 inst_12017 ( .A(net_11311), .Z(net_11865) );
NAND2_X2 inst_4647 ( .ZN(net_2343), .A1(net_2342), .A2(net_2341) );
CLKBUF_X2 inst_18758 ( .A(net_12433), .Z(net_18606) );
DFFR_X1 inst_7408 ( .D(net_5702), .CK(net_14042), .RN(x6501), .Q(x306) );
NAND2_X2 inst_4709 ( .ZN(net_4371), .A1(net_1802), .A2(net_1713) );
CLKBUF_X2 inst_10461 ( .A(net_10308), .Z(net_10309) );
CLKBUF_X2 inst_15436 ( .A(net_15283), .Z(net_15284) );
CLKBUF_X2 inst_10820 ( .A(net_10466), .Z(net_10668) );
DFFR_X2 inst_7060 ( .QN(net_6809), .D(net_4618), .CK(net_11844), .RN(x6501) );
OAI21_X2 inst_3130 ( .B2(net_2282), .ZN(net_2193), .A(net_2192), .B1(net_682) );
NOR2_X2 inst_3347 ( .ZN(net_5578), .A1(net_5440), .A2(net_5439) );
CLKBUF_X2 inst_9568 ( .A(net_9415), .Z(net_9416) );
CLKBUF_X2 inst_11446 ( .A(net_11293), .Z(net_11294) );
NAND2_X2 inst_4136 ( .ZN(net_5385), .A1(net_5219), .A2(net_5002) );
INV_X4 inst_5341 ( .ZN(net_2473), .A(net_1289) );
CLKBUF_X2 inst_12585 ( .A(net_12432), .Z(net_12433) );
CLKBUF_X2 inst_17573 ( .A(net_17420), .Z(net_17421) );
CLKBUF_X2 inst_9372 ( .A(net_9219), .Z(net_9220) );
CLKBUF_X2 inst_9653 ( .A(net_9500), .Z(net_9501) );
MUX2_X2 inst_4985 ( .A(net_9042), .Z(net_3941), .B(net_3533), .S(net_622) );
INV_X4 inst_5164 ( .ZN(net_3163), .A(net_3037) );
CLKBUF_X2 inst_9461 ( .A(net_9161), .Z(net_9309) );
CLKBUF_X2 inst_9736 ( .A(net_9304), .Z(net_9584) );
CLKBUF_X2 inst_15971 ( .A(net_15818), .Z(net_15819) );
SDFF_X2 inst_1655 ( .SI(net_7709), .Q(net_7709), .D(net_2659), .SE(net_2559), .CK(net_18538) );
CLKBUF_X2 inst_10720 ( .A(net_10567), .Z(net_10568) );
CLKBUF_X2 inst_15174 ( .A(net_15021), .Z(net_15022) );
DFFR_X1 inst_7415 ( .D(net_5725), .CK(net_13822), .RN(x6501), .Q(x9) );
CLKBUF_X2 inst_14165 ( .A(net_14012), .Z(net_14013) );
AOI221_X4 inst_8731 ( .B1(net_8884), .C1(net_8329), .B2(net_6252), .ZN(net_6221), .C2(net_4345), .A(net_4242) );
CLKBUF_X2 inst_16200 ( .A(net_9520), .Z(net_16048) );
CLKBUF_X2 inst_16594 ( .A(net_16441), .Z(net_16442) );
NAND2_X2 inst_4847 ( .A2(net_6820), .A1(net_2015), .ZN(net_1393) );
INV_X4 inst_6010 ( .A(net_6461), .ZN(net_3292) );
CLKBUF_X2 inst_16318 ( .A(net_12112), .Z(net_16166) );
CLKBUF_X2 inst_15733 ( .A(net_15580), .Z(net_15581) );
SDFF_X2 inst_1066 ( .D(net_7318), .SI(net_6494), .Q(net_6494), .SE(net_3071), .CK(net_12102) );
CLKBUF_X2 inst_9978 ( .A(net_9825), .Z(net_9826) );
AOI22_X2 inst_7977 ( .B1(net_7924), .A1(net_7822), .B2(net_6103), .A2(net_4398), .ZN(net_4153) );
CLKBUF_X2 inst_16542 ( .A(net_16389), .Z(net_16390) );
CLKBUF_X2 inst_10377 ( .A(net_10224), .Z(net_10225) );
CLKBUF_X2 inst_12122 ( .A(net_11969), .Z(net_11970) );
INV_X4 inst_5063 ( .ZN(net_5937), .A(net_5935) );
CLKBUF_X2 inst_15707 ( .A(net_12481), .Z(net_15555) );
NAND2_X2 inst_4608 ( .A2(net_6144), .ZN(net_2625), .A1(net_2624) );
SDFFR_X2 inst_2294 ( .SE(net_2260), .Q(net_329), .D(net_329), .CK(net_11519), .RN(x6501), .SI(x2693) );
CLKBUF_X2 inst_16909 ( .A(net_16756), .Z(net_16757) );
CLKBUF_X2 inst_14321 ( .A(net_14168), .Z(net_14169) );
CLKBUF_X2 inst_12495 ( .A(net_10366), .Z(net_12343) );
NAND2_X2 inst_4821 ( .ZN(net_1171), .A2(net_822), .A1(net_170) );
AOI222_X1 inst_8696 ( .C2(net_5832), .A2(net_5830), .B2(net_5824), .ZN(net_3202), .A1(net_2566), .B1(net_2131), .C1(x3156) );
NAND3_X2 inst_3931 ( .ZN(net_5531), .A1(net_5284), .A3(net_4792), .A2(net_4689) );
CLKBUF_X2 inst_12409 ( .A(net_12163), .Z(net_12257) );
CLKBUF_X2 inst_12682 ( .A(net_12529), .Z(net_12530) );
DFFR_X2 inst_7239 ( .QN(net_6393), .D(net_2226), .CK(net_15670), .RN(x6501) );
CLKBUF_X2 inst_13237 ( .A(net_9668), .Z(net_13085) );
CLKBUF_X2 inst_11590 ( .A(net_11437), .Z(net_11438) );
CLKBUF_X2 inst_10785 ( .A(net_9370), .Z(net_10633) );
CLKBUF_X2 inst_13098 ( .A(net_12868), .Z(net_12946) );
AOI221_X2 inst_8864 ( .C1(net_7212), .A(net_2528), .ZN(net_1728), .C2(net_1727), .B2(net_1622), .B1(net_602) );
XNOR2_X2 inst_158 ( .B(net_4884), .ZN(net_1938), .A(net_1849) );
CLKBUF_X2 inst_13529 ( .A(net_9791), .Z(net_13377) );
SDFF_X2 inst_507 ( .SI(net_8601), .Q(net_8601), .SE(net_3984), .D(net_3937), .CK(net_13051) );
NAND2_X2 inst_4289 ( .A1(net_6889), .A2(net_5247), .ZN(net_5171) );
CLKBUF_X2 inst_10566 ( .A(net_10413), .Z(net_10414) );
CLKBUF_X2 inst_14365 ( .A(net_14212), .Z(net_14213) );
SDFF_X2 inst_884 ( .Q(net_8563), .D(net_8563), .SI(net_3981), .SE(net_3878), .CK(net_10135) );
CLKBUF_X2 inst_12311 ( .A(net_12158), .Z(net_12159) );
SDFF_X2 inst_711 ( .SI(net_8639), .Q(net_8639), .D(net_3946), .SE(net_3885), .CK(net_11066) );
INV_X2 inst_6542 ( .A(net_6751), .ZN(net_3068) );
CLKBUF_X2 inst_14452 ( .A(net_11335), .Z(net_14300) );
CLKBUF_X2 inst_18847 ( .A(net_18694), .Z(net_18695) );
CLKBUF_X2 inst_14845 ( .A(net_12497), .Z(net_14693) );
CLKBUF_X2 inst_17559 ( .A(net_17406), .Z(net_17407) );
AOI22_X2 inst_8465 ( .B1(net_6738), .A1(net_6705), .B2(net_6202), .A2(net_3520), .ZN(net_3475) );
CLKBUF_X2 inst_11213 ( .A(net_11060), .Z(net_11061) );
CLKBUF_X2 inst_16725 ( .A(net_10811), .Z(net_16573) );
NAND2_X2 inst_4191 ( .ZN(net_5309), .A1(net_5065), .A2(net_5064) );
NAND2_X2 inst_4269 ( .A1(net_6916), .A2(net_5247), .ZN(net_5191) );
CLKBUF_X2 inst_14171 ( .A(net_14018), .Z(net_14019) );
CLKBUF_X2 inst_18581 ( .A(net_18428), .Z(net_18429) );
CLKBUF_X2 inst_18486 ( .A(net_15947), .Z(net_18334) );
AOI22_X2 inst_8559 ( .A1(net_2762), .ZN(net_2557), .B2(net_2556), .A2(net_2305), .B1(net_2123) );
CLKBUF_X2 inst_17936 ( .A(net_10072), .Z(net_17784) );
CLKBUF_X2 inst_15616 ( .A(net_15463), .Z(net_15464) );
CLKBUF_X2 inst_14534 ( .A(net_12971), .Z(net_14382) );
SDFFR_X2 inst_2263 ( .D(net_7380), .SE(net_2802), .SI(net_189), .Q(net_189), .CK(net_14974), .RN(x6501) );
INV_X4 inst_5608 ( .A(net_7503), .ZN(net_4459) );
NAND2_X2 inst_4796 ( .A1(net_2836), .ZN(net_2479), .A2(net_1256) );
NOR2_X2 inst_3549 ( .ZN(net_1441), .A2(net_1440), .A1(net_1065) );
NOR2_X2 inst_3501 ( .ZN(net_1863), .A1(net_1862), .A2(net_1861) );
CLKBUF_X2 inst_12602 ( .A(net_10704), .Z(net_12450) );
CLKBUF_X2 inst_10035 ( .A(net_9882), .Z(net_9883) );
CLKBUF_X2 inst_13029 ( .A(net_9354), .Z(net_12877) );
NAND2_X2 inst_4175 ( .ZN(net_5332), .A1(net_5193), .A2(net_4989) );
DFFR_X2 inst_7076 ( .QN(net_8295), .D(net_3970), .CK(net_11240), .RN(x6501) );
AOI22_X2 inst_8535 ( .B1(net_6592), .A1(net_6559), .A2(net_6257), .B2(net_6110), .ZN(net_3405) );
CLKBUF_X2 inst_9783 ( .A(net_9630), .Z(net_9631) );
CLKBUF_X2 inst_14217 ( .A(net_14064), .Z(net_14065) );
DFFS_X1 inst_6954 ( .D(net_3231), .CK(net_16332), .SN(x6501), .Q(x912) );
DFFR_X1 inst_7378 ( .D(net_5910), .CK(net_17192), .RN(x6501), .Q(x154) );
CLKBUF_X2 inst_9416 ( .A(net_9263), .Z(net_9264) );
NAND2_X2 inst_4397 ( .A1(net_7045), .A2(net_5162), .ZN(net_5060) );
OAI21_X2 inst_3102 ( .ZN(net_2579), .A(net_2577), .B2(net_2260), .B1(net_724) );
DFFR_X1 inst_7392 ( .QN(net_6299), .D(net_5855), .CK(net_16777), .RN(x6501) );
CLKBUF_X2 inst_10818 ( .A(net_9258), .Z(net_10666) );
CLKBUF_X2 inst_12847 ( .A(net_12694), .Z(net_12695) );
NAND4_X2 inst_3860 ( .A1(net_2829), .A4(net_2752), .A3(net_2493), .ZN(net_2454), .A2(net_1053) );
CLKBUF_X2 inst_12748 ( .A(net_12595), .Z(net_12596) );
SDFFS_X2 inst_2063 ( .SI(net_7393), .SE(net_2417), .Q(net_182), .D(net_182), .CK(net_17746), .SN(x6501) );
CLKBUF_X2 inst_14659 ( .A(net_9222), .Z(net_14507) );
CLKBUF_X2 inst_14917 ( .A(net_14764), .Z(net_14765) );
NAND2_X2 inst_4801 ( .A1(net_1522), .ZN(net_1373), .A2(net_1372) );
NAND4_X2 inst_3723 ( .ZN(net_4307), .A1(net_4178), .A2(net_4177), .A3(net_4176), .A4(net_4175) );
CLKBUF_X2 inst_15978 ( .A(net_15825), .Z(net_15826) );
CLKBUF_X2 inst_9346 ( .A(net_9109), .Z(net_9194) );
CLKBUF_X2 inst_12286 ( .A(net_12133), .Z(net_12134) );
CLKBUF_X2 inst_15282 ( .A(net_10911), .Z(net_15130) );
SDFF_X2 inst_2036 ( .SI(net_7913), .Q(net_7913), .D(net_2659), .SE(net_2461), .CK(net_15380) );
NAND3_X2 inst_3985 ( .ZN(net_1832), .A3(net_1556), .A2(net_967), .A1(net_935) );
INV_X4 inst_5386 ( .ZN(net_1335), .A(net_1178) );
CLKBUF_X2 inst_14350 ( .A(net_13282), .Z(net_14198) );
CLKBUF_X2 inst_9853 ( .A(net_9700), .Z(net_9701) );
CLKBUF_X2 inst_11107 ( .A(net_9947), .Z(net_10955) );
SDFF_X2 inst_868 ( .Q(net_8577), .D(net_8577), .SI(net_3956), .SE(net_3878), .CK(net_13233) );
SDFF_X2 inst_2049 ( .SI(net_7918), .Q(net_7918), .D(net_2584), .SE(net_2461), .CK(net_15561) );
AOI22_X2 inst_8187 ( .B1(net_8864), .A1(net_8309), .B2(net_6252), .A2(net_4345), .ZN(net_3845) );
CLKBUF_X2 inst_10747 ( .A(net_9504), .Z(net_10595) );
INV_X16 inst_6625 ( .ZN(net_4399), .A(net_3562) );
XNOR2_X2 inst_201 ( .B(net_6468), .ZN(net_1543), .A(net_1542) );
CLKBUF_X2 inst_11240 ( .A(net_11087), .Z(net_11088) );
NAND4_X2 inst_3627 ( .ZN(net_5599), .A2(net_5530), .A4(net_4864), .A1(net_4662), .A3(net_4531) );
XNOR2_X2 inst_304 ( .B(net_7367), .ZN(net_971), .A(net_970) );
SDFF_X2 inst_1084 ( .D(net_7338), .SI(net_6514), .Q(net_6514), .SE(net_3071), .CK(net_9470) );
NAND2_X2 inst_4157 ( .ZN(net_5357), .A1(net_5205), .A2(net_4995) );
INV_X4 inst_5793 ( .A(net_6364), .ZN(net_545) );
SDFF_X2 inst_1345 ( .SI(net_7273), .Q(net_7090), .D(net_7090), .SE(net_6278), .CK(net_14150) );
CLKBUF_X2 inst_10670 ( .A(net_10517), .Z(net_10518) );
CLKBUF_X2 inst_12823 ( .A(net_12670), .Z(net_12671) );
OAI222_X2 inst_2947 ( .C1(net_8214), .ZN(net_3891), .C2(net_3889), .A2(net_3888), .B2(net_3887), .A1(net_3600), .B1(net_693) );
CLKBUF_X2 inst_17650 ( .A(net_9646), .Z(net_17498) );
INV_X4 inst_5122 ( .ZN(net_5520), .A(net_4409) );
CLKBUF_X2 inst_12951 ( .A(net_12798), .Z(net_12799) );
CLKBUF_X2 inst_14225 ( .A(net_14072), .Z(net_14073) );
INV_X4 inst_5638 ( .A(net_7476), .ZN(net_3113) );
NOR2_X2 inst_3608 ( .ZN(net_1160), .A1(net_1093), .A2(net_845) );
DFFR_X2 inst_7306 ( .D(net_7631), .Q(net_7626), .CK(net_11213), .RN(x6501) );
CLKBUF_X2 inst_10724 ( .A(net_10213), .Z(net_10572) );
CLKBUF_X2 inst_15235 ( .A(net_15082), .Z(net_15083) );
SDFF_X2 inst_1016 ( .SI(net_7312), .Q(net_6653), .D(net_6653), .SE(net_3126), .CK(net_12026) );
CLKBUF_X2 inst_18195 ( .A(net_18042), .Z(net_18043) );
SDFF_X2 inst_848 ( .SI(net_8660), .Q(net_8660), .D(net_3940), .SE(net_3885), .CK(net_10321) );
CLKBUF_X2 inst_17480 ( .A(net_17327), .Z(net_17328) );
CLKBUF_X2 inst_13394 ( .A(net_13241), .Z(net_13242) );
SDFFR_X2 inst_2479 ( .Q(net_8973), .D(net_8973), .SI(net_4732), .SE(net_2562), .CK(net_14808), .RN(x6501) );
CLKBUF_X2 inst_14333 ( .A(net_14180), .Z(net_14181) );
CLKBUF_X2 inst_19153 ( .A(net_19000), .Z(net_19001) );
CLKBUF_X2 inst_17814 ( .A(net_17411), .Z(net_17662) );
SDFF_X2 inst_1554 ( .Q(net_7982), .D(net_7982), .SI(net_2708), .SE(net_2542), .CK(net_18273) );
CLKBUF_X2 inst_19162 ( .A(net_19009), .Z(net_19010) );
SDFF_X2 inst_1542 ( .Q(net_7997), .D(net_7997), .SI(net_2713), .SE(net_2542), .CK(net_16507) );
NAND2_X2 inst_4511 ( .A2(net_6207), .ZN(net_4368), .A1(net_4275) );
AOI22_X2 inst_7830 ( .B2(net_5535), .ZN(net_4691), .A2(net_4562), .A1(net_2701), .B1(net_444) );
AOI221_X2 inst_8849 ( .B1(net_8870), .C1(net_8315), .B2(net_6252), .ZN(net_6247), .C2(net_4345), .A(net_4258) );
CLKBUF_X2 inst_11580 ( .A(net_11427), .Z(net_11428) );
SDFF_X2 inst_644 ( .SI(net_8527), .Q(net_8527), .SE(net_3979), .D(net_3937), .CK(net_11080) );
CLKBUF_X2 inst_15946 ( .A(net_15793), .Z(net_15794) );
INV_X8 inst_5015 ( .ZN(net_5268), .A(net_4954) );
CLKBUF_X2 inst_19122 ( .A(net_12023), .Z(net_18970) );
CLKBUF_X2 inst_17229 ( .A(net_11932), .Z(net_17077) );
OR3_X2 inst_2806 ( .A3(net_3080), .ZN(net_2855), .A2(x12843), .A1(x12780) );
NAND3_X2 inst_4008 ( .A1(net_9014), .ZN(net_2531), .A2(net_1084), .A3(net_894) );
DFF_X1 inst_6736 ( .Q(net_6781), .D(net_5633), .CK(net_11430) );
INV_X2 inst_6449 ( .A(net_7560), .ZN(net_597) );
CLKBUF_X2 inst_10652 ( .A(net_9194), .Z(net_10500) );
CLKBUF_X2 inst_12229 ( .A(net_12076), .Z(net_12077) );
NAND2_X2 inst_4896 ( .A2(net_7386), .ZN(net_648), .A1(net_175) );
CLKBUF_X2 inst_14800 ( .A(net_10134), .Z(net_14648) );
SDFF_X2 inst_432 ( .Q(net_8742), .D(net_8742), .SE(net_3982), .SI(net_3943), .CK(net_13147) );
XNOR2_X2 inst_282 ( .ZN(net_1018), .B(net_939), .A(net_204) );
CLKBUF_X2 inst_16827 ( .A(net_9359), .Z(net_16675) );
CLKBUF_X2 inst_15829 ( .A(net_15676), .Z(net_15677) );
AOI21_X2 inst_8906 ( .B2(net_5871), .ZN(net_5753), .A(net_5752), .B1(net_2725) );
CLKBUF_X2 inst_11584 ( .A(net_11431), .Z(net_11432) );
AOI22_X2 inst_8428 ( .B1(net_6531), .A1(net_6498), .A2(net_6137), .B2(net_6104), .ZN(net_3513) );
CLKBUF_X2 inst_9605 ( .A(net_9452), .Z(net_9453) );
CLKBUF_X2 inst_12533 ( .A(net_11445), .Z(net_12381) );
OAI21_X2 inst_3171 ( .ZN(net_1244), .B1(net_1243), .B2(net_955), .A(net_899) );
NOR3_X2 inst_3266 ( .A1(net_2967), .ZN(net_2839), .A3(net_2424), .A2(net_2307) );
AOI221_X4 inst_8725 ( .B1(net_8838), .C1(net_8357), .C2(net_6265), .B2(net_6253), .ZN(net_4340), .A(net_4252) );
CLKBUF_X2 inst_14060 ( .A(net_11038), .Z(net_13908) );
CLKBUF_X2 inst_14910 ( .A(net_14757), .Z(net_14758) );
CLKBUF_X2 inst_12479 ( .A(net_12326), .Z(net_12327) );
CLKBUF_X2 inst_18681 ( .A(net_18528), .Z(net_18529) );
CLKBUF_X2 inst_18106 ( .A(net_17953), .Z(net_17954) );
AOI22_X2 inst_7887 ( .B1(net_8999), .A2(net_5609), .B2(net_5456), .ZN(net_4544), .A1(net_378) );
CLKBUF_X2 inst_10296 ( .A(net_10143), .Z(net_10144) );
SDFF_X2 inst_774 ( .Q(net_8785), .D(net_8785), .SI(net_3981), .SE(net_3879), .CK(net_12950) );
SDFFR_X2 inst_2292 ( .SE(net_5582), .D(net_2635), .CK(net_14198), .RN(x6501), .SI(x105), .Q(x105) );
CLKBUF_X2 inst_16418 ( .A(net_16265), .Z(net_16266) );
CLKBUF_X2 inst_14826 ( .A(net_10018), .Z(net_14674) );
CLKBUF_X2 inst_16871 ( .A(net_16718), .Z(net_16719) );
INV_X4 inst_5300 ( .A(net_2043), .ZN(net_1686) );
SDFFR_X1 inst_2766 ( .QN(net_7579), .D(net_3958), .SE(net_3144), .SI(net_626), .CK(net_10954), .RN(x6501) );
CLKBUF_X2 inst_12340 ( .A(net_12187), .Z(net_12188) );
NAND2_X2 inst_4326 ( .A1(net_7140), .A2(net_5166), .ZN(net_5131) );
AOI22_X2 inst_7938 ( .B1(net_8157), .A1(net_7715), .B2(net_6101), .A2(net_6095), .ZN(net_6002) );
CLKBUF_X2 inst_13985 ( .A(net_13832), .Z(net_13833) );
CLKBUF_X2 inst_18663 ( .A(net_18510), .Z(net_18511) );
CLKBUF_X2 inst_18382 ( .A(net_12123), .Z(net_18230) );
XNOR2_X2 inst_127 ( .ZN(net_2866), .B(net_2807), .A(net_2806) );
CLKBUF_X2 inst_14754 ( .A(net_11606), .Z(net_14602) );
CLKBUF_X2 inst_17535 ( .A(net_17382), .Z(net_17383) );
CLKBUF_X2 inst_11279 ( .A(net_9637), .Z(net_11127) );
CLKBUF_X2 inst_10657 ( .A(net_10504), .Z(net_10505) );
CLKBUF_X2 inst_14562 ( .A(net_14409), .Z(net_14410) );
XNOR2_X2 inst_122 ( .ZN(net_2930), .A(net_2811), .B(net_890) );
SDFF_X2 inst_1268 ( .Q(net_7813), .D(net_7813), .SE(net_2730), .SI(net_2658), .CK(net_15554) );
OAI21_X2 inst_3029 ( .B2(net_4971), .ZN(net_4937), .A(net_4789), .B1(net_756) );
CLKBUF_X2 inst_14270 ( .A(net_14117), .Z(net_14118) );
AOI21_X2 inst_8944 ( .B2(net_5784), .ZN(net_5604), .A(net_5600), .B1(net_2673) );
CLKBUF_X2 inst_15053 ( .A(net_14900), .Z(net_14901) );
CLKBUF_X2 inst_9740 ( .A(net_9587), .Z(net_9588) );
INV_X2 inst_6281 ( .ZN(net_4220), .A(net_3933) );
DFFR_X1 inst_7540 ( .QN(net_7630), .D(net_2021), .CK(net_11186), .RN(x6501) );
CLKBUF_X2 inst_17657 ( .A(net_17504), .Z(net_17505) );
NAND3_X2 inst_3912 ( .ZN(net_5626), .A1(net_5555), .A3(net_5489), .A2(net_5346) );
CLKBUF_X2 inst_10077 ( .A(net_9221), .Z(net_9925) );
AOI22_X2 inst_8499 ( .B1(net_6614), .A1(net_6581), .A2(net_6257), .B2(net_6110), .ZN(net_3441) );
SDFFR_X2 inst_2306 ( .SE(net_2260), .Q(net_334), .D(net_334), .CK(net_11481), .RN(x6501), .SI(x2451) );
AND2_X2 inst_9191 ( .ZN(net_1849), .A2(net_1677), .A1(net_754) );
SDFF_X2 inst_1646 ( .SI(net_7724), .Q(net_7724), .D(net_2718), .SE(net_2559), .CK(net_14914) );
CLKBUF_X2 inst_14008 ( .A(net_13855), .Z(net_13856) );
CLKBUF_X2 inst_14468 ( .A(net_14315), .Z(net_14316) );
CLKBUF_X2 inst_15361 ( .A(net_12191), .Z(net_15209) );
DFF_X1 inst_6748 ( .Q(net_6759), .D(net_5617), .CK(net_10499) );
INV_X4 inst_5773 ( .A(net_7597), .ZN(net_1016) );
DFFR_X1 inst_7547 ( .Q(net_8266), .D(net_3550), .CK(net_18506), .RN(x6501) );
CLKBUF_X2 inst_17167 ( .A(net_17014), .Z(net_17015) );
INV_X2 inst_6294 ( .ZN(net_4204), .A(net_3913) );
DFF_X1 inst_6741 ( .Q(net_6785), .D(net_5628), .CK(net_11425) );
CLKBUF_X2 inst_13664 ( .A(net_10524), .Z(net_13512) );
CLKBUF_X2 inst_18536 ( .A(net_18383), .Z(net_18384) );
INV_X4 inst_5550 ( .ZN(net_1092), .A(net_894) );
SDFF_X2 inst_1102 ( .D(net_7331), .SI(net_6540), .Q(net_6540), .SE(net_3086), .CK(net_9421) );
INV_X2 inst_6368 ( .ZN(net_2310), .A(net_1719) );
CLKBUF_X2 inst_13329 ( .A(net_13176), .Z(net_13177) );
SDFF_X2 inst_702 ( .Q(net_8426), .D(net_8426), .SI(net_3958), .SE(net_3934), .CK(net_10000) );
INV_X4 inst_5860 ( .A(net_6360), .ZN(net_535) );
CLKBUF_X2 inst_12448 ( .A(net_11357), .Z(net_12296) );
CLKBUF_X2 inst_18668 ( .A(net_13821), .Z(net_18516) );
CLKBUF_X2 inst_15192 ( .A(net_15039), .Z(net_15040) );
CLKBUF_X2 inst_9297 ( .A(net_9144), .Z(net_9145) );
CLKBUF_X2 inst_9980 ( .A(net_9117), .Z(net_9828) );
CLKBUF_X2 inst_12233 ( .A(net_12080), .Z(net_12081) );
CLKBUF_X2 inst_13912 ( .A(net_13363), .Z(net_13760) );
AND3_X2 inst_9049 ( .ZN(net_1881), .A1(net_1704), .A3(net_1703), .A2(net_1521) );
CLKBUF_X2 inst_18533 ( .A(net_18315), .Z(net_18381) );
CLKBUF_X2 inst_12365 ( .A(net_10148), .Z(net_12213) );
OAI22_X2 inst_2928 ( .A1(net_3162), .B1(net_2931), .ZN(net_2838), .A2(net_2642), .B2(net_1711) );
CLKBUF_X2 inst_13335 ( .A(net_11587), .Z(net_13183) );
SDFF_X2 inst_400 ( .SI(net_8312), .Q(net_8312), .SE(net_3978), .D(net_3973), .CK(net_12357) );
NAND4_X2 inst_3813 ( .ZN(net_3613), .A1(net_3435), .A2(net_3434), .A3(net_3433), .A4(net_3432) );
OAI21_X2 inst_2991 ( .ZN(net_5903), .B2(net_5902), .A(net_5820), .B1(net_696) );
AOI21_X2 inst_8895 ( .B2(net_5871), .ZN(net_5791), .A(net_5790), .B1(x291) );
NOR2_X2 inst_3513 ( .A2(net_3023), .ZN(net_1774), .A1(net_1189) );
INV_X2 inst_6309 ( .ZN(net_3895), .A(net_3592) );
CLKBUF_X2 inst_16196 ( .A(net_16043), .Z(net_16044) );
XNOR2_X2 inst_261 ( .A(net_2744), .B(net_2688), .ZN(net_1183) );
CLKBUF_X2 inst_12418 ( .A(net_9841), .Z(net_12266) );
XNOR2_X2 inst_268 ( .A(net_6304), .B(net_2687), .ZN(net_1069) );
SDFF_X2 inst_1518 ( .Q(net_7886), .D(net_7886), .SI(net_2574), .SE(net_2543), .CK(net_15602) );
AOI22_X2 inst_8198 ( .B1(net_8718), .A1(net_8496), .B2(net_4350), .A2(net_4349), .ZN(net_3838) );
CLKBUF_X2 inst_10985 ( .A(net_10832), .Z(net_10833) );
AOI222_X4 inst_8586 ( .C1(net_7441), .A2(net_6266), .ZN(net_4416), .B2(net_4365), .C2(net_4364), .B1(net_4314), .A1(x13654) );
AND2_X2 inst_9199 ( .ZN(net_1582), .A1(net_1308), .A2(net_1307) );
CLKBUF_X2 inst_18313 ( .A(net_12142), .Z(net_18161) );
CLKBUF_X2 inst_12264 ( .A(net_12111), .Z(net_12112) );
CLKBUF_X2 inst_18092 ( .A(net_16809), .Z(net_17940) );
DFFR_X2 inst_7245 ( .QN(net_7399), .D(net_2052), .CK(net_17875), .RN(x6501) );
CLKBUF_X2 inst_14118 ( .A(net_13965), .Z(net_13966) );
NOR2_X2 inst_3509 ( .A2(net_2400), .A1(net_2397), .ZN(net_2113) );
CLKBUF_X2 inst_13936 ( .A(net_13783), .Z(net_13784) );
CLKBUF_X2 inst_17758 ( .A(net_11684), .Z(net_17606) );
AOI22_X2 inst_7971 ( .B1(net_8025), .A1(net_7991), .B2(net_6102), .A2(net_6097), .ZN(net_4158) );
CLKBUF_X2 inst_10746 ( .A(net_10416), .Z(net_10594) );
CLKBUF_X2 inst_11511 ( .A(net_9459), .Z(net_11359) );
INV_X2 inst_6348 ( .ZN(net_2404), .A(net_2403) );
OAI21_X2 inst_3097 ( .ZN(net_2771), .A(net_2765), .B2(net_1984), .B1(net_633) );
AOI22_X2 inst_8357 ( .B1(net_8813), .A1(net_8554), .A2(net_3861), .B2(net_3860), .ZN(net_3691) );
CLKBUF_X2 inst_9229 ( .A(net_9076), .Z(net_9077) );
CLKBUF_X2 inst_9625 ( .A(net_9472), .Z(net_9473) );
SDFF_X2 inst_502 ( .SI(net_8629), .Q(net_8629), .SE(net_3984), .D(net_3948), .CK(net_13428) );
CLKBUF_X2 inst_13976 ( .A(net_10023), .Z(net_13824) );
AOI221_X2 inst_8745 ( .B1(net_7197), .C2(net_6448), .ZN(net_5656), .B2(net_5655), .C1(net_5654), .A(net_5528) );
CLKBUF_X2 inst_18212 ( .A(net_16556), .Z(net_18060) );
CLKBUF_X2 inst_17966 ( .A(net_17813), .Z(net_17814) );
CLKBUF_X2 inst_14771 ( .A(net_11979), .Z(net_14619) );
NAND4_X2 inst_3645 ( .ZN(net_4916), .A3(net_4675), .A2(net_4549), .A4(net_4548), .A1(net_4464) );
SDFF_X2 inst_1598 ( .Q(net_8132), .D(net_8132), .SI(net_2718), .SE(net_2541), .CK(net_18787) );
CLKBUF_X2 inst_15724 ( .A(net_15228), .Z(net_15572) );
CLKBUF_X2 inst_17040 ( .A(net_14427), .Z(net_16888) );
CLKBUF_X2 inst_17098 ( .A(net_16945), .Z(net_16946) );
CLKBUF_X2 inst_10167 ( .A(net_10014), .Z(net_10015) );
CLKBUF_X2 inst_15670 ( .A(net_15517), .Z(net_15518) );
AOI22_X2 inst_7880 ( .A2(net_5538), .ZN(net_4552), .B1(net_4551), .B2(net_4388), .A1(net_422) );
OAI21_X2 inst_3152 ( .B2(net_1984), .ZN(net_1982), .A(net_1974), .B1(net_699) );
CLKBUF_X2 inst_15073 ( .A(net_12842), .Z(net_14921) );
NAND2_X2 inst_4161 ( .ZN(net_5352), .A1(net_5095), .A2(net_5094) );
CLKBUF_X2 inst_18166 ( .A(net_18013), .Z(net_18014) );
CLKBUF_X2 inst_11678 ( .A(net_11525), .Z(net_11526) );
CLKBUF_X2 inst_10117 ( .A(net_9964), .Z(net_9965) );
INV_X4 inst_5869 ( .A(net_8932), .ZN(net_2596) );
OAI211_X2 inst_3196 ( .C2(net_8893), .ZN(net_3154), .B(net_3153), .C1(net_3000), .A(net_1423) );
CLKBUF_X2 inst_14603 ( .A(net_14450), .Z(net_14451) );
INV_X2 inst_6525 ( .A(net_6805), .ZN(net_527) );
CLKBUF_X2 inst_15452 ( .A(net_15299), .Z(net_15300) );
CLKBUF_X2 inst_18252 ( .A(net_18099), .Z(net_18100) );
NAND2_X4 inst_4025 ( .A2(net_6084), .A1(net_6083), .ZN(net_3221) );
XNOR2_X2 inst_322 ( .A(net_7379), .B(net_1023), .ZN(net_938) );
NOR2_X2 inst_3516 ( .A2(net_1773), .ZN(net_1772), .A1(net_1521) );
CLKBUF_X2 inst_10070 ( .A(net_9461), .Z(net_9918) );
NAND2_X2 inst_4200 ( .ZN(net_5297), .A1(net_5056), .A2(net_5055) );
NAND3_X2 inst_3902 ( .ZN(net_5636), .A1(net_5565), .A3(net_5499), .A2(net_5386) );
INV_X2 inst_6191 ( .ZN(net_5736), .A(net_5735) );
CLKBUF_X2 inst_10858 ( .A(net_10705), .Z(net_10706) );
CLKBUF_X2 inst_10647 ( .A(net_9494), .Z(net_10495) );
INV_X2 inst_6243 ( .ZN(net_4863), .A(net_4766) );
DFFS_X2 inst_6908 ( .QN(net_6805), .D(net_6802), .CK(net_9625), .SN(x6501) );
AOI22_X2 inst_8302 ( .B1(net_8769), .A1(net_8399), .A2(net_3867), .B2(net_3866), .ZN(net_3742) );
INV_X2 inst_6289 ( .ZN(net_4210), .A(net_3918) );
SDFFR_X2 inst_2315 ( .SE(net_2260), .Q(net_358), .D(net_358), .CK(net_11514), .RN(x6501), .SI(x2006) );
CLKBUF_X2 inst_12662 ( .A(net_12509), .Z(net_12510) );
SDFF_X2 inst_962 ( .SI(net_7311), .Q(net_6718), .D(net_6718), .SE(net_3124), .CK(net_12128) );
INV_X2 inst_6350 ( .ZN(net_2312), .A(net_2220) );
CLKBUF_X2 inst_18789 ( .A(net_17363), .Z(net_18637) );
CLKBUF_X2 inst_11489 ( .A(net_10210), .Z(net_11337) );
CLKBUF_X2 inst_9673 ( .A(net_9267), .Z(net_9521) );
AOI22_X2 inst_7955 ( .B1(net_8057), .A1(net_7853), .B2(net_6107), .A2(net_4400), .ZN(net_4172) );
CLKBUF_X2 inst_17395 ( .A(net_15838), .Z(net_17243) );
CLKBUF_X2 inst_14044 ( .A(net_13891), .Z(net_13892) );
CLKBUF_X2 inst_19119 ( .A(net_18966), .Z(net_18967) );
CLKBUF_X2 inst_9308 ( .A(net_9109), .Z(net_9156) );
CLKBUF_X2 inst_11876 ( .A(net_11723), .Z(net_11724) );
SDFF_X2 inst_350 ( .SI(net_8466), .Q(net_8466), .SE(net_3983), .D(net_3956), .CK(net_13300) );
CLKBUF_X2 inst_11322 ( .A(net_11169), .Z(net_11170) );
CLKBUF_X2 inst_10403 ( .A(net_10250), .Z(net_10251) );
CLKBUF_X2 inst_14437 ( .A(net_14284), .Z(net_14285) );
INV_X4 inst_5104 ( .ZN(net_5673), .A(net_5603) );
CLKBUF_X2 inst_16853 ( .A(net_11474), .Z(net_16701) );
CLKBUF_X2 inst_18275 ( .A(net_18122), .Z(net_18123) );
CLKBUF_X2 inst_12851 ( .A(net_12698), .Z(net_12699) );
AOI22_X2 inst_8518 ( .B1(net_6684), .A1(net_6651), .A2(net_6213), .B2(net_6138), .ZN(net_3422) );
CLKBUF_X2 inst_11901 ( .A(net_11748), .Z(net_11749) );
DFFR_X1 inst_7506 ( .D(net_1706), .CK(net_16381), .RN(x6501), .Q(x963) );
SDFF_X2 inst_1452 ( .SI(net_7269), .Q(net_7086), .D(net_7086), .SE(net_6278), .CK(net_16853) );
CLKBUF_X2 inst_11867 ( .A(net_11714), .Z(net_11715) );
CLKBUF_X2 inst_13740 ( .A(net_13587), .Z(net_13588) );
INV_X2 inst_6549 ( .A(net_6362), .ZN(net_2125) );
CLKBUF_X2 inst_16743 ( .A(net_16590), .Z(net_16591) );
CLKBUF_X2 inst_18176 ( .A(net_18023), .Z(net_18024) );
CLKBUF_X2 inst_12967 ( .A(net_12814), .Z(net_12815) );
SDFF_X2 inst_1396 ( .SI(net_7725), .Q(net_7725), .D(net_2713), .SE(net_2559), .CK(net_16511) );
AOI21_X2 inst_8901 ( .B2(net_5871), .ZN(net_5779), .A(net_5752), .B1(x170) );
CLKBUF_X2 inst_15768 ( .A(net_15615), .Z(net_15616) );
CLKBUF_X2 inst_15311 ( .A(net_15158), .Z(net_15159) );
CLKBUF_X2 inst_16774 ( .A(net_16621), .Z(net_16622) );
OAI21_X2 inst_3003 ( .B2(net_5902), .ZN(net_5890), .A(net_5822), .B1(net_766) );
INV_X4 inst_5579 ( .A(net_6370), .ZN(net_780) );
CLKBUF_X2 inst_12169 ( .A(net_11355), .Z(net_12017) );
CLKBUF_X2 inst_16978 ( .A(net_16825), .Z(net_16826) );
CLKBUF_X2 inst_16641 ( .A(net_16488), .Z(net_16489) );
SDFFR_X2 inst_2185 ( .SI(net_7636), .Q(net_7636), .SE(net_3022), .D(net_1168), .CK(net_18914), .RN(x6501) );
AOI22_X2 inst_8550 ( .B2(net_4889), .A1(net_4803), .ZN(net_3333), .B1(net_3332), .A2(net_3199) );
AND2_X2 inst_9165 ( .A2(net_6105), .ZN(net_2662), .A1(net_2661) );
CLKBUF_X2 inst_13134 ( .A(net_12981), .Z(net_12982) );
NAND2_X4 inst_4050 ( .ZN(net_6251), .A1(net_2027), .A2(net_1561) );
CLKBUF_X2 inst_16604 ( .A(net_16451), .Z(net_16452) );
SDFFR_X2 inst_2370 ( .SE(net_2260), .Q(net_325), .D(net_325), .CK(net_10438), .RN(x6501), .SI(x2908) );
NAND3_X2 inst_3882 ( .ZN(net_5889), .A3(net_5777), .A1(net_4964), .A2(net_4785) );
CLKBUF_X2 inst_14069 ( .A(net_9589), .Z(net_13917) );
CLKBUF_X2 inst_16868 ( .A(net_16715), .Z(net_16716) );
OR3_X2 inst_2811 ( .A3(net_7618), .A2(net_2021), .ZN(net_1564), .A1(net_1563) );
CLKBUF_X2 inst_17597 ( .A(net_17444), .Z(net_17445) );
XNOR2_X2 inst_137 ( .ZN(net_2537), .A(net_2535), .B(net_1940) );
NAND2_X2 inst_4615 ( .A2(net_6144), .ZN(net_2611), .A1(net_2610) );
INV_X4 inst_6120 ( .A(net_9005), .ZN(net_483) );
CLKBUF_X2 inst_18067 ( .A(net_16630), .Z(net_17915) );
DFFS_X2 inst_6889 ( .Q(net_8964), .D(net_2890), .CK(net_14822), .SN(x6501) );
SDFFR_X2 inst_2567 ( .QN(net_6362), .SE(net_2147), .D(net_2125), .SI(net_1943), .CK(net_14655), .RN(x6501) );
CLKBUF_X2 inst_11384 ( .A(net_11231), .Z(net_11232) );
OAI211_X2 inst_3206 ( .C2(net_5036), .ZN(net_2637), .B(net_2155), .A(net_1514), .C1(net_1163) );
CLKBUF_X2 inst_11742 ( .A(net_11589), .Z(net_11590) );
AOI222_X2 inst_8591 ( .B2(net_6451), .B1(net_5654), .C2(net_5595), .A2(net_4881), .ZN(net_4707), .C1(net_333), .A1(net_251) );
CLKBUF_X2 inst_17576 ( .A(net_17423), .Z(net_17424) );
NAND2_X4 inst_4046 ( .ZN(net_2558), .A2(net_2267), .A1(net_2261) );
CLKBUF_X2 inst_10245 ( .A(net_10092), .Z(net_10093) );
DFFR_X2 inst_7179 ( .QN(net_6395), .D(net_2488), .CK(net_15680), .RN(x6501) );
CLKBUF_X2 inst_11752 ( .A(net_11599), .Z(net_11600) );
AOI22_X2 inst_8112 ( .B1(net_8013), .A1(net_7979), .B2(net_6102), .A2(net_6097), .ZN(net_5992) );
SDFF_X2 inst_1897 ( .D(net_7275), .SI(net_6852), .Q(net_6852), .SE(net_6282), .CK(net_14609) );
AOI22_X2 inst_8511 ( .B1(net_6616), .A1(net_6583), .A2(net_6257), .B2(net_6110), .ZN(net_3429) );
CLKBUF_X2 inst_18634 ( .A(net_18481), .Z(net_18482) );
CLKBUF_X2 inst_10615 ( .A(net_10462), .Z(net_10463) );
CLKBUF_X2 inst_11810 ( .A(net_10822), .Z(net_11658) );
OAI21_X2 inst_3159 ( .B2(net_2048), .ZN(net_1969), .A(net_1968), .B1(net_1862) );
CLKBUF_X2 inst_15587 ( .A(net_15434), .Z(net_15435) );
CLKBUF_X2 inst_15786 ( .A(net_15633), .Z(net_15634) );
SDFF_X2 inst_1569 ( .Q(net_8034), .D(net_8034), .SI(net_2717), .SE(net_2545), .CK(net_14406) );
DFFR_X2 inst_7130 ( .QN(net_7602), .D(net_3077), .CK(net_9778), .RN(x6501) );
CLKBUF_X2 inst_11722 ( .A(net_11569), .Z(net_11570) );
CLKBUF_X2 inst_12990 ( .A(net_12837), .Z(net_12838) );
SDFF_X2 inst_1772 ( .SI(net_8075), .Q(net_8075), .D(net_2716), .SE(net_2508), .CK(net_17060) );
DFFR_X2 inst_7080 ( .Q(net_7649), .D(net_3896), .CK(net_12688), .RN(x6501) );
DFFR_X2 inst_7314 ( .Q(net_394), .D(net_392), .CK(net_13859), .RN(x6501) );
CLKBUF_X2 inst_13565 ( .A(net_13412), .Z(net_13413) );
CLKBUF_X2 inst_13725 ( .A(net_13572), .Z(net_13573) );
CLKBUF_X2 inst_14738 ( .A(net_14585), .Z(net_14586) );
SDFFR_X2 inst_2143 ( .SI(net_7182), .Q(net_7182), .D(net_6433), .SE(net_4362), .CK(net_16428), .RN(x6501) );
SDFF_X2 inst_1291 ( .Q(net_7824), .D(net_7824), .SE(net_2730), .SI(net_2590), .CK(net_18415) );
CLKBUF_X2 inst_14233 ( .A(net_14080), .Z(net_14081) );
SDFF_X2 inst_359 ( .SI(net_8305), .Q(net_8305), .SE(net_3978), .D(net_3937), .CK(net_12483) );
AOI22_X2 inst_8239 ( .B1(net_8742), .A1(net_8372), .A2(net_3867), .B2(net_3866), .ZN(net_3798) );
CLKBUF_X2 inst_18030 ( .A(net_17877), .Z(net_17878) );
CLKBUF_X2 inst_12382 ( .A(net_10556), .Z(net_12230) );
SDFF_X2 inst_1962 ( .D(net_7283), .SI(net_6900), .Q(net_6900), .SE(net_6284), .CK(net_18979) );
NAND2_X2 inst_4757 ( .ZN(net_2450), .A2(net_2012), .A1(net_1670) );
CLKBUF_X2 inst_13037 ( .A(net_11293), .Z(net_12885) );
CLKBUF_X2 inst_13582 ( .A(net_13429), .Z(net_13430) );
CLKBUF_X2 inst_10492 ( .A(net_9360), .Z(net_10340) );
CLKBUF_X2 inst_11551 ( .A(net_11398), .Z(net_11399) );
CLKBUF_X2 inst_15334 ( .A(net_15181), .Z(net_15182) );
INV_X4 inst_5283 ( .ZN(net_1628), .A(net_1528) );
CLKBUF_X2 inst_12925 ( .A(net_12772), .Z(net_12773) );
CLKBUF_X2 inst_15635 ( .A(net_15482), .Z(net_15483) );
INV_X2 inst_6174 ( .ZN(net_5931), .A(net_5923) );
AOI22_X2 inst_8168 ( .B1(net_8751), .A1(net_8381), .ZN(net_3868), .A2(net_3867), .B2(net_3866) );
XNOR2_X2 inst_194 ( .ZN(net_1551), .B(net_1199), .A(net_1197) );
AOI22_X2 inst_8421 ( .B1(net_6728), .A1(net_6695), .B2(net_6202), .ZN(net_3521), .A2(net_3520) );
NOR2_X2 inst_3453 ( .A1(net_3023), .ZN(net_2928), .A2(net_2867) );
CLKBUF_X2 inst_15594 ( .A(net_15441), .Z(net_15442) );
CLKBUF_X2 inst_14181 ( .A(net_11588), .Z(net_14029) );
INV_X4 inst_6136 ( .A(net_7208), .ZN(net_1787) );
AOI221_X4 inst_8714 ( .C1(net_7939), .B1(net_7837), .C2(net_6103), .ZN(net_6051), .B2(net_4398), .A(net_4286) );
CLKBUF_X2 inst_11317 ( .A(net_11164), .Z(net_11165) );
SDFF_X2 inst_442 ( .Q(net_8771), .D(net_8771), .SE(net_3982), .SI(net_3940), .CK(net_10290) );
SDFFR_X2 inst_2507 ( .Q(net_9001), .D(net_9001), .SI(net_4743), .SE(net_2562), .CK(net_16401), .RN(x6501) );
AOI22_X2 inst_8338 ( .B1(net_8847), .A1(net_8366), .A2(net_6265), .B2(net_6253), .ZN(net_3709) );
CLKBUF_X2 inst_9337 ( .A(net_9184), .Z(net_9185) );
SDFFR_X2 inst_2245 ( .SE(net_2802), .D(net_2785), .SI(net_190), .Q(net_190), .CK(net_14992), .RN(x6501) );
CLKBUF_X2 inst_14751 ( .A(net_11950), .Z(net_14599) );
INV_X4 inst_5237 ( .ZN(net_2265), .A(net_2192) );
CLKBUF_X2 inst_12620 ( .A(net_12467), .Z(net_12468) );
CLKBUF_X2 inst_15467 ( .A(net_11469), .Z(net_15315) );
INV_X4 inst_6097 ( .A(net_7600), .ZN(net_1186) );
NAND2_X2 inst_4298 ( .A1(net_7051), .A2(net_5162), .ZN(net_5159) );
CLKBUF_X2 inst_11242 ( .A(net_9899), .Z(net_11090) );
CLKBUF_X2 inst_14593 ( .A(net_14440), .Z(net_14441) );
SDFF_X2 inst_1249 ( .SI(net_7694), .Q(net_7694), .D(net_2717), .SE(net_2714), .CK(net_14189) );
DFFR_X2 inst_7212 ( .D(net_2374), .QN(net_207), .CK(net_17792), .RN(x6501) );
NAND2_X2 inst_4099 ( .ZN(net_5435), .A2(net_5244), .A1(net_5156) );
CLKBUF_X2 inst_15815 ( .A(net_14965), .Z(net_15663) );
NAND2_X2 inst_4740 ( .ZN(net_2575), .A2(net_1586), .A1(net_978) );
INV_X4 inst_5403 ( .ZN(net_1144), .A(net_879) );
INV_X4 inst_5967 ( .A(net_7568), .ZN(net_515) );
SDFF_X2 inst_1318 ( .SI(net_7703), .Q(net_7703), .SE(net_2714), .D(net_2703), .CK(net_14027) );
DFFS_X2 inst_6894 ( .D(net_2761), .QN(net_186), .CK(net_14997), .SN(x6501) );
DFFR_X2 inst_7219 ( .D(net_2364), .QN(net_210), .CK(net_17883), .RN(x6501) );
CLKBUF_X2 inst_16970 ( .A(net_16817), .Z(net_16818) );
CLKBUF_X2 inst_18444 ( .A(net_18291), .Z(net_18292) );
SDFF_X2 inst_1070 ( .D(net_7323), .SI(net_6532), .Q(net_6532), .SE(net_3086), .CK(net_11354) );
NAND2_X2 inst_4584 ( .ZN(net_2910), .A1(net_2909), .A2(net_2908) );
SDFFR_X2 inst_2454 ( .D(net_4884), .SE(net_2685), .SI(net_408), .Q(net_408), .CK(net_13930), .RN(x6501) );
CLKBUF_X2 inst_12037 ( .A(net_11884), .Z(net_11885) );
NOR2_X2 inst_3601 ( .ZN(net_1274), .A1(net_1273), .A2(net_841) );
CLKBUF_X2 inst_12255 ( .A(net_9166), .Z(net_12103) );
CLKBUF_X2 inst_14612 ( .A(net_14459), .Z(net_14460) );
CLKBUF_X2 inst_9693 ( .A(net_9227), .Z(net_9541) );
NAND2_X2 inst_4536 ( .ZN(net_3375), .A1(net_3374), .A2(net_3373) );
CLKBUF_X2 inst_18840 ( .A(net_18687), .Z(net_18688) );
INV_X4 inst_5601 ( .A(net_7405), .ZN(net_751) );
CLKBUF_X2 inst_11854 ( .A(net_11339), .Z(net_11702) );
DFF_X1 inst_6763 ( .Q(net_7543), .D(net_4609), .CK(net_9731) );
SDFF_X2 inst_1673 ( .SI(net_7742), .Q(net_7742), .D(net_2709), .SE(net_2560), .CK(net_15751) );
INV_X4 inst_5745 ( .A(net_8941), .ZN(net_6219) );
CLKBUF_X2 inst_15163 ( .A(net_15010), .Z(net_15011) );
CLKBUF_X2 inst_18832 ( .A(net_11321), .Z(net_18680) );
CLKBUF_X2 inst_14373 ( .A(net_14220), .Z(net_14221) );
SDFF_X2 inst_1153 ( .SI(net_7335), .Q(net_6610), .D(net_6610), .SE(net_3069), .CK(net_9749) );
NAND4_X2 inst_3823 ( .ZN(net_3603), .A1(net_3395), .A2(net_3394), .A3(net_3393), .A4(net_3392) );
AOI22_X2 inst_7959 ( .B1(net_8024), .A1(net_7990), .B2(net_6102), .A2(net_6097), .ZN(net_6036) );
DFFR_X2 inst_7325 ( .D(net_7642), .QN(net_7639), .CK(net_15646), .RN(x6501) );
CLKBUF_X2 inst_10905 ( .A(net_10752), .Z(net_10753) );
SDFF_X2 inst_391 ( .Q(net_8841), .D(net_8841), .SI(net_3975), .SE(net_3964), .CK(net_12559) );
CLKBUF_X2 inst_18272 ( .A(net_18119), .Z(net_18120) );
CLKBUF_X2 inst_19165 ( .A(net_19012), .Z(net_19013) );
NAND2_X2 inst_4107 ( .ZN(net_5424), .A1(net_5149), .A2(net_5148) );
CLKBUF_X2 inst_15020 ( .A(net_13094), .Z(net_14868) );
CLKBUF_X2 inst_18014 ( .A(net_17861), .Z(net_17862) );
CLKBUF_X2 inst_17939 ( .A(net_17786), .Z(net_17787) );
CLKBUF_X2 inst_14092 ( .A(net_9118), .Z(net_13940) );
AOI22_X2 inst_8035 ( .B1(net_8203), .A1(net_7693), .B2(net_6099), .A2(net_4399), .ZN(net_4103) );
CLKBUF_X2 inst_10896 ( .A(net_10743), .Z(net_10744) );
INV_X4 inst_6074 ( .A(net_5963), .ZN(x2981) );
CLKBUF_X2 inst_17702 ( .A(net_17549), .Z(net_17550) );
CLKBUF_X2 inst_17045 ( .A(net_16892), .Z(net_16893) );
AOI22_X2 inst_8403 ( .B1(net_8823), .A1(net_8342), .A2(net_6265), .B2(net_6253), .ZN(net_3649) );
SDFF_X2 inst_1799 ( .D(net_7285), .SI(net_6982), .Q(net_6982), .SE(net_6283), .CK(net_19008) );
NAND2_X2 inst_4442 ( .A1(net_6879), .A2(net_5016), .ZN(net_4985) );
CLKBUF_X2 inst_15129 ( .A(net_10811), .Z(net_14977) );
DFFR_X1 inst_7385 ( .D(net_5860), .CK(net_11497), .RN(x6501), .Q(x3604) );
CLKBUF_X2 inst_9326 ( .A(net_9173), .Z(net_9174) );
CLKBUF_X2 inst_17954 ( .A(net_17801), .Z(net_17802) );
NOR2_X2 inst_3458 ( .A1(net_3023), .ZN(net_2823), .A2(net_2746) );
SDFF_X2 inst_1313 ( .SI(net_7701), .Q(net_7701), .D(net_2716), .SE(net_2714), .CK(net_16872) );
NAND2_X2 inst_4694 ( .A1(net_7559), .ZN(net_1903), .A2(net_1729) );
AOI22_X2 inst_8098 ( .A1(net_7973), .B1(net_7803), .A2(net_6092), .B2(net_6091), .ZN(net_4049) );
CLKBUF_X2 inst_11104 ( .A(net_9405), .Z(net_10952) );
CLKBUF_X2 inst_14572 ( .A(net_10843), .Z(net_14420) );
AOI222_X1 inst_8632 ( .A2(net_6266), .ZN(net_4366), .B2(net_4365), .C2(net_4364), .B1(net_3991), .C1(net_3990), .A1(x13733) );
CLKBUF_X2 inst_16192 ( .A(net_16039), .Z(net_16040) );
OR2_X2 inst_2886 ( .A2(net_2077), .ZN(net_1869), .A1(net_1797) );
NAND2_X2 inst_4116 ( .ZN(net_5412), .A1(net_5140), .A2(net_5139) );
CLKBUF_X2 inst_15146 ( .A(net_14993), .Z(net_14994) );
CLKBUF_X2 inst_14851 ( .A(net_14557), .Z(net_14699) );
INV_X2 inst_6523 ( .ZN(net_530), .A(x13208) );
INV_X4 inst_5150 ( .ZN(net_3189), .A(net_3164) );
CLKBUF_X2 inst_9613 ( .A(net_9460), .Z(net_9461) );
CLKBUF_X2 inst_13747 ( .A(net_13594), .Z(net_13595) );
CLKBUF_X2 inst_10978 ( .A(net_10825), .Z(net_10826) );
SDFFS_X2 inst_2081 ( .SI(net_7377), .SE(net_2794), .Q(net_166), .D(net_166), .CK(net_17733), .SN(x6501) );
SDFFR_X1 inst_2773 ( .D(net_7382), .Q(net_7279), .SI(net_1950), .SE(net_1327), .CK(net_14659), .RN(x6501) );
CLKBUF_X2 inst_13199 ( .A(net_13046), .Z(net_13047) );
NOR3_X2 inst_3261 ( .ZN(net_3232), .A1(net_3193), .A3(net_1037), .A2(net_875) );
AOI221_X4 inst_8717 ( .B1(net_8714), .C1(net_8492), .ZN(net_4352), .B2(net_4350), .C2(net_4349), .A(net_4266) );
CLKBUF_X2 inst_16570 ( .A(net_16417), .Z(net_16418) );
CLKBUF_X2 inst_13606 ( .A(net_13174), .Z(net_13454) );
CLKBUF_X2 inst_15796 ( .A(net_12455), .Z(net_15644) );
SDFF_X2 inst_1211 ( .Q(net_7965), .D(net_7965), .SE(net_2755), .SI(net_2749), .CK(net_13802) );
SDFF_X2 inst_1192 ( .D(net_7310), .SI(net_6552), .Q(net_6552), .SE(net_3086), .CK(net_11852) );
SDFF_X2 inst_682 ( .Q(net_8692), .D(net_8692), .SI(net_3954), .SE(net_3935), .CK(net_13247) );
XNOR2_X2 inst_238 ( .ZN(net_1239), .B(net_874), .A(net_515) );
CLKBUF_X2 inst_12394 ( .A(net_11269), .Z(net_12242) );
CLKBUF_X2 inst_16012 ( .A(net_15859), .Z(net_15860) );
CLKBUF_X2 inst_16338 ( .A(net_16185), .Z(net_16186) );
NOR2_X4 inst_3333 ( .A2(net_6200), .ZN(net_5832), .A1(net_2986) );
CLKBUF_X2 inst_15908 ( .A(net_15755), .Z(net_15756) );
CLKBUF_X2 inst_10021 ( .A(net_9868), .Z(net_9869) );
OAI21_X2 inst_3109 ( .B1(net_2731), .ZN(net_2481), .A(net_2480), .B2(net_2479) );
CLKBUF_X2 inst_10046 ( .A(net_9893), .Z(net_9894) );
CLKBUF_X2 inst_18448 ( .A(net_18295), .Z(net_18296) );
SDFFR_X2 inst_2240 ( .Q(net_7459), .D(net_7459), .SE(net_2863), .CK(net_10617), .SI(x13514), .RN(x6501) );
CLKBUF_X2 inst_14995 ( .A(net_14842), .Z(net_14843) );
SDFF_X2 inst_1210 ( .Q(net_7970), .D(net_7970), .SE(net_2755), .SI(net_2715), .CK(net_14308) );
CLKBUF_X2 inst_11680 ( .A(net_11527), .Z(net_11528) );
INV_X4 inst_6090 ( .A(net_7561), .ZN(net_3145) );
CLKBUF_X2 inst_12759 ( .A(net_12606), .Z(net_12607) );
CLKBUF_X2 inst_14674 ( .A(net_14521), .Z(net_14522) );
CLKBUF_X2 inst_17804 ( .A(net_14755), .Z(net_17652) );
SDFFR_X2 inst_2437 ( .D(net_2671), .SE(net_2313), .SI(net_458), .Q(net_458), .CK(net_13830), .RN(x6501) );
CLKBUF_X2 inst_15154 ( .A(net_14361), .Z(net_15002) );
CLKBUF_X2 inst_18553 ( .A(net_18400), .Z(net_18401) );
NAND2_X2 inst_4521 ( .ZN(net_3575), .A1(net_3574), .A2(net_3573) );
AOI22_X2 inst_8324 ( .B1(net_8845), .A1(net_8364), .A2(net_6265), .B2(net_6253), .ZN(net_3722) );
SDFF_X2 inst_1981 ( .D(net_7295), .SI(net_6912), .Q(net_6912), .SE(net_6284), .CK(net_15390) );
INV_X2 inst_6324 ( .ZN(net_3339), .A(net_3281) );
INV_X4 inst_5960 ( .A(net_9012), .ZN(net_1084) );
CLKBUF_X2 inst_18190 ( .A(net_15784), .Z(net_18038) );
CLKBUF_X2 inst_15122 ( .A(net_14969), .Z(net_14970) );
CLKBUF_X2 inst_17022 ( .A(net_16869), .Z(net_16870) );
AOI22_X2 inst_8309 ( .B1(net_8585), .A1(net_8474), .A2(net_6263), .B2(net_6262), .ZN(net_3736) );
NAND4_X2 inst_3775 ( .ZN(net_4246), .A1(net_3737), .A2(net_3736), .A3(net_3735), .A4(net_3734) );
CLKBUF_X2 inst_16266 ( .A(net_16113), .Z(net_16114) );
CLKBUF_X2 inst_13762 ( .A(net_13609), .Z(net_13610) );
SDFFR_X2 inst_2472 ( .SE(net_2678), .D(net_2569), .SI(net_437), .Q(net_437), .CK(net_14541), .RN(x6501) );
CLKBUF_X2 inst_14900 ( .A(net_13960), .Z(net_14748) );
CLKBUF_X2 inst_11239 ( .A(net_11086), .Z(net_11087) );
AOI22_X2 inst_8293 ( .B1(net_8768), .A1(net_8398), .A2(net_3867), .B2(net_3866), .ZN(net_3749) );
SDFF_X2 inst_872 ( .Q(net_8583), .D(net_8583), .SI(net_3941), .SE(net_3878), .CK(net_12498) );
INV_X16 inst_6641 ( .ZN(net_3861), .A(net_3317) );
CLKBUF_X2 inst_16795 ( .A(net_16642), .Z(net_16643) );
CLKBUF_X2 inst_11479 ( .A(net_11326), .Z(net_11327) );
CLKBUF_X2 inst_14821 ( .A(net_14668), .Z(net_14669) );
CLKBUF_X2 inst_9210 ( .A(x12768), .Z(net_9058) );
INV_X4 inst_5234 ( .A(net_2649), .ZN(net_2198) );
CLKBUF_X2 inst_12579 ( .A(net_12426), .Z(net_12427) );
CLKBUF_X2 inst_14907 ( .A(net_14754), .Z(net_14755) );
SDFF_X2 inst_1667 ( .SI(net_7764), .Q(net_7764), .D(net_2710), .SE(net_2560), .CK(net_14401) );
CLKBUF_X2 inst_15375 ( .A(net_15222), .Z(net_15223) );
CLKBUF_X2 inst_17985 ( .A(net_15043), .Z(net_17833) );
SDFF_X2 inst_462 ( .SI(net_8465), .Q(net_8465), .SE(net_3983), .D(net_3957), .CK(net_13277) );
CLKBUF_X2 inst_15339 ( .A(net_15186), .Z(net_15187) );
CLKBUF_X2 inst_10261 ( .A(net_10108), .Z(net_10109) );
INV_X4 inst_5572 ( .A(net_6819), .ZN(net_2015) );
CLKBUF_X2 inst_9398 ( .A(net_9245), .Z(net_9246) );
CLKBUF_X2 inst_10579 ( .A(net_10426), .Z(net_10427) );
DFFR_X2 inst_7223 ( .QN(net_7666), .D(net_2258), .CK(net_14574), .RN(x6501) );
CLKBUF_X2 inst_18975 ( .A(net_14687), .Z(net_18823) );
CLKBUF_X2 inst_18641 ( .A(net_18488), .Z(net_18489) );
CLKBUF_X2 inst_13381 ( .A(net_13228), .Z(net_13229) );
HA_X1 inst_6661 ( .S(net_3583), .CO(net_3582), .A(net_3581), .B(net_3270) );
CLKBUF_X2 inst_18693 ( .A(net_18540), .Z(net_18541) );
CLKBUF_X2 inst_10389 ( .A(net_9494), .Z(net_10237) );
NAND2_X1 inst_4909 ( .A1(net_2043), .ZN(net_1610), .A2(net_383) );
DFFR_X2 inst_7114 ( .QN(net_7610), .D(net_3058), .CK(net_9811), .RN(x6501) );
DFF_X1 inst_6836 ( .Q(net_6455), .D(net_3612), .CK(net_15155) );
SDFF_X2 inst_1914 ( .D(net_7283), .SI(net_7020), .Q(net_7020), .SE(net_6277), .CK(net_16172) );
SDFF_X2 inst_1975 ( .D(net_7267), .SI(net_7004), .Q(net_7004), .SE(net_6277), .CK(net_16795) );
INV_X2 inst_6219 ( .ZN(net_5491), .A(net_5353) );
CLKBUF_X2 inst_14702 ( .A(net_14549), .Z(net_14550) );
CLKBUF_X2 inst_15855 ( .A(net_11214), .Z(net_15703) );
INV_X16 inst_6647 ( .ZN(net_6099), .A(net_3564) );
NAND2_X2 inst_4806 ( .A1(net_8953), .A2(net_2466), .ZN(net_1310) );
CLKBUF_X2 inst_9728 ( .A(net_9575), .Z(net_9576) );
CLKBUF_X2 inst_9585 ( .A(net_9338), .Z(net_9433) );
AOI22_X2 inst_8117 ( .B1(net_8149), .A1(net_7707), .B2(net_6101), .A2(net_6095), .ZN(net_4031) );
CLKBUF_X2 inst_12362 ( .A(net_12209), .Z(net_12210) );
CLKBUF_X2 inst_17944 ( .A(net_17791), .Z(net_17792) );
CLKBUF_X2 inst_17155 ( .A(net_17002), .Z(net_17003) );
CLKBUF_X2 inst_11893 ( .A(net_11740), .Z(net_11741) );
OAI21_X2 inst_3017 ( .ZN(net_5045), .B2(net_5044), .A(net_4892), .B1(net_1312) );
INV_X2 inst_6389 ( .A(net_3161), .ZN(net_1276) );
CLKBUF_X2 inst_17693 ( .A(net_12179), .Z(net_17541) );
SDFF_X2 inst_845 ( .SI(net_8657), .Q(net_8657), .D(net_3941), .SE(net_3885), .CK(net_12864) );
NOR2_X2 inst_3554 ( .A2(net_3320), .A1(net_3318), .ZN(net_1370) );
SDFF_X2 inst_1367 ( .Q(net_8211), .D(net_8211), .SI(net_2716), .SE(net_2561), .CK(net_14290) );
CLKBUF_X2 inst_17613 ( .A(net_9619), .Z(net_17461) );
CLKBUF_X2 inst_17289 ( .A(net_17136), .Z(net_17137) );
CLKBUF_X2 inst_10980 ( .A(net_9236), .Z(net_10828) );
AND2_X2 inst_9175 ( .A2(net_6188), .ZN(net_2392), .A1(net_2391) );
CLKBUF_X2 inst_16911 ( .A(net_12342), .Z(net_16759) );
CLKBUF_X2 inst_10898 ( .A(net_10745), .Z(net_10746) );
NAND4_X2 inst_3687 ( .A4(net_6242), .A1(net_6241), .ZN(net_4450), .A2(net_3844), .A3(net_3843) );
CLKBUF_X2 inst_15426 ( .A(net_13746), .Z(net_15274) );
CLKBUF_X2 inst_10837 ( .A(net_10684), .Z(net_10685) );
AOI22_X2 inst_8434 ( .B1(net_6665), .A1(net_6632), .A2(net_6213), .B2(net_6138), .ZN(net_3507) );
CLKBUF_X2 inst_17676 ( .A(net_13200), .Z(net_17524) );
CLKBUF_X2 inst_10103 ( .A(net_9257), .Z(net_9951) );
OAI21_X2 inst_3053 ( .B2(net_8234), .B1(net_4850), .ZN(net_4758), .A(net_2611) );
AOI22_X2 inst_7829 ( .A2(net_5657), .B2(net_5463), .ZN(net_4692), .A1(net_2641), .B1(net_435) );
CLKBUF_X2 inst_10409 ( .A(net_10256), .Z(net_10257) );
NAND2_X2 inst_4810 ( .A2(net_2556), .ZN(net_1285), .A1(net_1284) );
CLKBUF_X2 inst_9962 ( .A(net_9809), .Z(net_9810) );
CLKBUF_X2 inst_10708 ( .A(net_10555), .Z(net_10556) );
CLKBUF_X2 inst_17202 ( .A(net_16467), .Z(net_17050) );
OAI21_X2 inst_3103 ( .ZN(net_2578), .A(net_2577), .B2(net_2260), .B1(net_629) );
CLKBUF_X2 inst_16075 ( .A(net_15922), .Z(net_15923) );
CLKBUF_X2 inst_11985 ( .A(net_11832), .Z(net_11833) );
NOR3_X2 inst_3304 ( .A2(net_2206), .A1(net_1740), .A3(net_1739), .ZN(net_1738) );
DFFR_X1 inst_7520 ( .Q(net_6417), .D(net_1102), .CK(net_9672), .RN(x6501) );
CLKBUF_X2 inst_16045 ( .A(net_15892), .Z(net_15893) );
AOI22_X2 inst_7762 ( .B1(net_6962), .A1(net_6922), .A2(net_5443), .B2(net_5442), .ZN(net_5358) );
INV_X4 inst_5384 ( .ZN(net_1517), .A(net_1103) );
CLKBUF_X2 inst_17275 ( .A(net_17122), .Z(net_17123) );
CLKBUF_X2 inst_16766 ( .A(net_16613), .Z(net_16614) );
NAND2_X2 inst_4723 ( .A1(net_7375), .ZN(net_1979), .A2(net_1783) );
NAND4_X2 inst_3655 ( .A4(net_6004), .A1(net_6003), .ZN(net_4610), .A2(net_4162), .A3(net_4161) );
DFFR_X1 inst_7532 ( .Q(net_7657), .D(net_919), .CK(net_12711), .RN(x6501) );
CLKBUF_X2 inst_12145 ( .A(net_9159), .Z(net_11993) );
HA_X1 inst_6692 ( .S(net_2920), .CO(net_2919), .B(net_2563), .A(x3258) );
INV_X2 inst_6617 ( .ZN(net_6211), .A(net_6209) );
SDFF_X2 inst_1888 ( .D(net_7266), .SI(net_6963), .Q(net_6963), .SE(net_6283), .CK(net_14337) );
OR2_X4 inst_2843 ( .ZN(net_2187), .A1(net_2156), .A2(net_1923) );
SDFF_X2 inst_1763 ( .D(net_7285), .SI(net_6942), .Q(net_6942), .SE(net_6281), .CK(net_19021) );
NOR2_X2 inst_3379 ( .ZN(net_5546), .A1(net_5309), .A2(net_5308) );
CLKBUF_X2 inst_13071 ( .A(net_12382), .Z(net_12919) );
CLKBUF_X2 inst_16061 ( .A(net_13803), .Z(net_15909) );
CLKBUF_X2 inst_18473 ( .A(net_18320), .Z(net_18321) );
DFFR_X2 inst_7190 ( .QN(net_8958), .D(net_2451), .CK(net_15068), .RN(x6501) );
CLKBUF_X2 inst_13685 ( .A(net_13532), .Z(net_13533) );
SDFF_X2 inst_1094 ( .D(net_7320), .SI(net_6496), .Q(net_6496), .SE(net_3071), .CK(net_12086) );
CLKBUF_X2 inst_14309 ( .A(net_14156), .Z(net_14157) );
NAND2_X2 inst_4145 ( .ZN(net_5373), .A1(net_5213), .A2(net_4999) );
CLKBUF_X2 inst_19179 ( .A(net_19026), .Z(net_19027) );
NAND2_X2 inst_4590 ( .A2(net_2881), .ZN(net_2880), .A1(net_1268) );
NAND4_X2 inst_3680 ( .A4(net_6032), .A1(net_6031), .ZN(net_4585), .A2(net_4010), .A3(net_4009) );
INV_X2 inst_6376 ( .A(net_2084), .ZN(net_1368) );
DFFR_X2 inst_7168 ( .QN(net_8903), .D(net_2581), .CK(net_16299), .RN(x6501) );
SDFF_X2 inst_1699 ( .SI(net_7722), .Q(net_7722), .D(net_2590), .SE(net_2559), .CK(net_15969) );
NAND2_X2 inst_4878 ( .ZN(net_1411), .A2(net_800), .A1(net_168) );
CLKBUF_X2 inst_12685 ( .A(net_11424), .Z(net_12533) );
XOR2_X2 inst_50 ( .B(net_3128), .Z(net_1005), .A(net_1004) );
CLKBUF_X2 inst_18906 ( .A(net_9076), .Z(net_18754) );
CLKBUF_X2 inst_16324 ( .A(net_16171), .Z(net_16172) );
SDFFR_X2 inst_2589 ( .QN(net_7257), .D(net_2760), .SI(net_1947), .SE(net_1379), .CK(net_18112), .RN(x6501) );
CLKBUF_X2 inst_11762 ( .A(net_11433), .Z(net_11610) );
CLKBUF_X2 inst_10626 ( .A(net_10473), .Z(net_10474) );
CLKBUF_X2 inst_16849 ( .A(net_16696), .Z(net_16697) );
AOI222_X1 inst_8699 ( .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_2970), .B1(net_2969), .C1(net_2968), .A2(net_2300) );
SDFF_X2 inst_1650 ( .SI(net_7732), .Q(net_7732), .D(net_2715), .SE(net_2559), .CK(net_14262) );
CLKBUF_X2 inst_18074 ( .A(net_17921), .Z(net_17922) );
CLKBUF_X2 inst_19098 ( .A(net_18945), .Z(net_18946) );
NAND2_X2 inst_4439 ( .A1(net_6876), .A2(net_5016), .ZN(net_4988) );
DFFR_X1 inst_7469 ( .QN(net_7439), .D(net_4270), .CK(net_12852), .RN(x6501) );
AOI22_X2 inst_8250 ( .B1(net_8873), .A1(net_8318), .B2(net_6252), .A2(net_4345), .ZN(net_3786) );
OR2_X2 inst_2872 ( .A1(net_4905), .A2(net_4834), .ZN(net_4641) );
AOI222_X1 inst_8683 ( .B1(net_6482), .A2(net_3296), .B2(net_3295), .C2(net_3294), .ZN(net_3289), .A1(net_3284), .C1(net_980) );
CLKBUF_X2 inst_18702 ( .A(net_16883), .Z(net_18550) );
NOR2_X2 inst_3380 ( .ZN(net_5545), .A1(net_5305), .A2(net_5304) );
CLKBUF_X2 inst_16887 ( .A(net_16734), .Z(net_16735) );
SDFF_X2 inst_804 ( .SI(net_8492), .Q(net_8492), .D(net_3960), .SE(net_3884), .CK(net_13094) );
CLKBUF_X2 inst_16147 ( .A(net_15994), .Z(net_15995) );
CLKBUF_X2 inst_15965 ( .A(net_11099), .Z(net_15813) );
NOR3_X2 inst_3290 ( .A3(net_2849), .ZN(net_2203), .A1(net_1996), .A2(net_1377) );
AOI221_X2 inst_8824 ( .C1(net_8156), .B1(net_7714), .C2(net_6101), .B2(net_6095), .ZN(net_5997), .A(net_4309) );
XOR2_X2 inst_13 ( .Z(net_1510), .A(net_1509), .B(net_1171) );
SDFFR_X2 inst_2584 ( .QN(net_7255), .SI(net_1953), .SE(net_1379), .D(net_1330), .CK(net_18113), .RN(x6501) );
CLKBUF_X2 inst_14527 ( .A(net_14374), .Z(net_14375) );
SDFFR_X1 inst_2755 ( .QN(net_7562), .D(net_3943), .SE(net_3144), .SI(net_3138), .CK(net_10960), .RN(x6501) );
AND2_X4 inst_9101 ( .ZN(net_2542), .A2(net_2267), .A1(net_2263) );
CLKBUF_X2 inst_9393 ( .A(net_9240), .Z(net_9241) );
CLKBUF_X2 inst_17443 ( .A(net_17290), .Z(net_17291) );
SDFF_X2 inst_1819 ( .D(net_7265), .SI(net_6842), .Q(net_6842), .SE(net_6282), .CK(net_14354) );
CLKBUF_X2 inst_14718 ( .A(net_12995), .Z(net_14566) );
CLKBUF_X2 inst_17080 ( .A(net_16927), .Z(net_16928) );
SDFF_X2 inst_453 ( .SI(net_8445), .Q(net_8445), .SE(net_3983), .D(net_3961), .CK(net_13210) );
SDFF_X2 inst_493 ( .SI(net_8618), .Q(net_8618), .SE(net_3984), .D(net_3954), .CK(net_12629) );
XOR2_X2 inst_23 ( .Z(net_1384), .B(net_1383), .A(net_706) );
SDFF_X2 inst_1822 ( .D(net_7284), .SI(net_6861), .Q(net_6861), .SE(net_6282), .CK(net_16197) );
NAND4_X2 inst_3790 ( .ZN(net_4231), .A1(net_3639), .A2(net_3638), .A3(net_3637), .A4(net_3636) );
CLKBUF_X2 inst_18765 ( .A(net_18612), .Z(net_18613) );
CLKBUF_X2 inst_12551 ( .A(net_11838), .Z(net_12399) );
CLKBUF_X2 inst_17282 ( .A(net_17030), .Z(net_17130) );
HA_X1 inst_6701 ( .CO(net_6136), .A(net_2968), .S(net_2300), .B(net_2038) );
CLKBUF_X2 inst_15574 ( .A(net_12679), .Z(net_15422) );
CLKBUF_X2 inst_10340 ( .A(net_10069), .Z(net_10188) );
CLKBUF_X2 inst_14798 ( .A(net_14645), .Z(net_14646) );
SDFF_X2 inst_812 ( .SI(net_8502), .Q(net_8502), .D(net_3957), .SE(net_3884), .CK(net_12332) );
CLKBUF_X2 inst_10347 ( .A(net_9797), .Z(net_10195) );
CLKBUF_X2 inst_15535 ( .A(net_15382), .Z(net_15383) );
XNOR2_X2 inst_179 ( .B(net_6380), .ZN(net_1699), .A(net_1599) );
CLKBUF_X2 inst_15603 ( .A(net_10003), .Z(net_15451) );
SDFF_X2 inst_1730 ( .Q(net_7989), .D(net_7989), .SI(net_2720), .SE(net_2542), .CK(net_15240) );
INV_X4 inst_5698 ( .A(net_6372), .ZN(net_571) );
NAND4_X2 inst_3799 ( .ZN(net_3627), .A2(net_3491), .A1(net_3490), .A3(net_3489), .A4(net_3488) );
XOR2_X1 inst_76 ( .Z(net_3279), .A(net_3165), .B(x2355) );
NAND4_X2 inst_3734 ( .ZN(net_4296), .A1(net_4112), .A2(net_4111), .A3(net_4110), .A4(net_4109) );
XNOR2_X2 inst_172 ( .B(net_2397), .ZN(net_1793), .A(net_1792) );
DFF_X1 inst_6769 ( .Q(net_7548), .D(net_4603), .CK(net_12773) );
CLKBUF_X2 inst_11228 ( .A(net_11075), .Z(net_11076) );
CLKBUF_X2 inst_16870 ( .A(net_9726), .Z(net_16718) );
XNOR2_X2 inst_277 ( .A(net_3550), .ZN(net_1031), .B(net_1020) );
NAND2_X2 inst_4366 ( .A1(net_7112), .A2(net_5164), .ZN(net_5091) );
XOR2_X1 inst_83 ( .B(net_3205), .Z(net_3017), .A(net_2870) );
AOI22_X2 inst_7787 ( .A2(net_6187), .ZN(net_4828), .B2(net_4555), .B1(net_2000), .A1(net_206) );
NAND2_X2 inst_4186 ( .ZN(net_5316), .A2(net_5186), .A1(net_5069) );
INV_X4 inst_5566 ( .A(net_1106), .ZN(net_601) );
AOI22_X2 inst_7946 ( .A1(net_7954), .B1(net_7784), .A2(net_6092), .B2(net_6091), .ZN(net_4180) );
NOR2_X2 inst_3386 ( .ZN(net_4686), .A1(net_4685), .A2(net_4684) );
CLKBUF_X2 inst_13673 ( .A(net_13520), .Z(net_13521) );
XNOR2_X2 inst_140 ( .ZN(net_2535), .A(net_2108), .B(net_2107) );
AOI22_X2 inst_7990 ( .B1(net_8130), .A1(net_7892), .A2(net_6098), .B2(net_4190), .ZN(net_4142) );
CLKBUF_X2 inst_16880 ( .A(net_16727), .Z(net_16728) );
OR2_X4 inst_2824 ( .A2(net_6205), .ZN(net_4559), .A1(net_1103) );
INV_X4 inst_5945 ( .A(net_6457), .ZN(net_2949) );
NOR2_X2 inst_3594 ( .ZN(net_1282), .A1(net_1084), .A2(net_894) );
AOI22_X2 inst_8155 ( .B1(net_8019), .A1(net_7985), .B2(net_6102), .A2(net_6097), .ZN(net_3997) );
OAI21_X2 inst_3124 ( .B2(net_2299), .ZN(net_2258), .A(net_2253), .B1(net_673) );
AOI22_X2 inst_7993 ( .B1(net_8198), .A1(net_7688), .B2(net_6099), .A2(net_4399), .ZN(net_4139) );
OAI221_X2 inst_2952 ( .C2(net_6456), .B2(net_6133), .ZN(net_4951), .C1(net_4950), .A(net_4828), .B1(net_1413) );
CLKBUF_X2 inst_11896 ( .A(net_11743), .Z(net_11744) );
CLKBUF_X2 inst_14990 ( .A(net_12794), .Z(net_14838) );
CLKBUF_X2 inst_17621 ( .A(net_17468), .Z(net_17469) );
XNOR2_X2 inst_174 ( .ZN(net_1789), .A(net_1788), .B(net_1461) );
CLKBUF_X2 inst_11558 ( .A(net_11405), .Z(net_11406) );
CLKBUF_X2 inst_17313 ( .A(net_17160), .Z(net_17161) );
CLKBUF_X2 inst_16462 ( .A(net_16309), .Z(net_16310) );
AOI222_X1 inst_8658 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3908), .B1(net_2923), .C1(net_2921), .A1(x13797) );
AOI21_X2 inst_8942 ( .A(net_5783), .ZN(net_5715), .B2(net_5519), .B1(net_5464) );
CLKBUF_X2 inst_12293 ( .A(net_12140), .Z(net_12141) );
XOR2_X2 inst_5 ( .Z(net_3091), .A(net_2919), .B(x3207) );
SDFFR_X2 inst_2105 ( .SE(net_5876), .Q(net_306), .D(net_306), .SI(net_257), .CK(net_14721), .RN(x6501) );
CLKBUF_X2 inst_11186 ( .A(net_11033), .Z(net_11034) );
CLKBUF_X2 inst_17718 ( .A(net_14541), .Z(net_17566) );
CLKBUF_X2 inst_17778 ( .A(net_17625), .Z(net_17626) );
SDFF_X2 inst_729 ( .SI(net_8343), .Q(net_8343), .D(net_3946), .SE(net_3880), .CK(net_10718) );
INV_X2 inst_6567 ( .A(net_8270), .ZN(net_488) );
SDFFR_X2 inst_2157 ( .Q(net_8276), .D(net_8276), .SI(net_8272), .SE(net_2996), .CK(net_18430), .RN(x6501) );
INV_X2 inst_6506 ( .A(net_6379), .ZN(net_2041) );
CLKBUF_X2 inst_10891 ( .A(net_9727), .Z(net_10739) );
SDFFR_X1 inst_2783 ( .D(net_7380), .Q(net_7277), .SI(net_1943), .SE(net_1327), .CK(net_14658), .RN(x6501) );
NAND2_X2 inst_4553 ( .ZN(net_3527), .A1(net_3359), .A2(net_3301) );
SDFF_X2 inst_604 ( .SI(net_8398), .Q(net_8398), .SE(net_3969), .D(net_3941), .CK(net_13414) );
INV_X4 inst_5804 ( .A(net_7601), .ZN(net_846) );
AOI211_X2 inst_9004 ( .A(net_7616), .ZN(net_5751), .C1(net_5691), .C2(net_5597), .B(net_5453) );
DFFR_X2 inst_7085 ( .Q(net_7653), .D(net_3886), .CK(net_10453), .RN(x6501) );
DFFR_X1 inst_7539 ( .Q(net_6480), .D(net_1542), .CK(net_11734), .RN(x6501) );
CLKBUF_X2 inst_13872 ( .A(net_13719), .Z(net_13720) );
NAND2_X2 inst_4057 ( .ZN(net_5918), .A2(net_5838), .A1(net_5588) );
SDFF_X2 inst_1179 ( .SI(net_7338), .Q(net_6613), .D(net_6613), .SE(net_3069), .CK(net_9440) );
XNOR2_X2 inst_292 ( .ZN(net_1000), .A(net_999), .B(net_975) );
NAND4_X2 inst_3650 ( .A4(net_5998), .A1(net_5997), .ZN(net_4615), .A2(net_4193), .A3(net_4192) );
CLKBUF_X2 inst_11661 ( .A(net_11508), .Z(net_11509) );
SDFF_X2 inst_2012 ( .SI(net_7777), .Q(net_7777), .D(net_2659), .SE(net_2459), .CK(net_18022) );
CLKBUF_X2 inst_11350 ( .A(net_11197), .Z(net_11198) );
CLKBUF_X2 inst_10900 ( .A(net_10747), .Z(net_10748) );
CLKBUF_X2 inst_16768 ( .A(net_15673), .Z(net_16616) );
INV_X2 inst_6605 ( .A(net_6164), .ZN(net_6163) );
SDFF_X2 inst_839 ( .SI(net_8631), .Q(net_8631), .D(net_3943), .SE(net_3885), .CK(net_13328) );
CLKBUF_X2 inst_16296 ( .A(net_16143), .Z(net_16144) );
XNOR2_X2 inst_240 ( .A(net_6837), .ZN(net_1222), .B(net_1221) );
INV_X4 inst_5455 ( .A(net_939), .ZN(net_854) );
NAND3_X2 inst_3966 ( .ZN(net_2470), .A1(net_2402), .A2(net_2401), .A3(net_1891) );
DFFR_X1 inst_7501 ( .Q(net_7263), .D(net_1879), .CK(net_14792), .RN(x6501) );
CLKBUF_X2 inst_13681 ( .A(net_13528), .Z(net_13529) );
XOR2_X1 inst_99 ( .B(net_3032), .A(net_2949), .Z(net_1215) );
INV_X16 inst_6634 ( .ZN(net_3863), .A(net_3365) );
CLKBUF_X2 inst_9997 ( .A(net_9844), .Z(net_9845) );
CLKBUF_X2 inst_13210 ( .A(net_13057), .Z(net_13058) );
CLKBUF_X2 inst_13152 ( .A(net_12999), .Z(net_13000) );
NAND2_X2 inst_4384 ( .A1(net_7118), .A2(net_5164), .ZN(net_5073) );
CLKBUF_X2 inst_11050 ( .A(net_10593), .Z(net_10898) );
SDFF_X2 inst_2059 ( .SI(net_7937), .Q(net_7937), .D(net_2660), .SE(net_2461), .CK(net_16957) );
CLKBUF_X2 inst_13851 ( .A(net_13698), .Z(net_13699) );
DFFR_X2 inst_7023 ( .QN(net_6302), .D(net_5696), .CK(net_16933), .RN(x6501) );
CLKBUF_X2 inst_9445 ( .A(net_9180), .Z(net_9293) );
CLKBUF_X2 inst_9473 ( .A(net_9320), .Z(net_9321) );
XNOR2_X2 inst_311 ( .ZN(net_960), .A(net_959), .B(net_958) );
CLKBUF_X2 inst_9656 ( .A(net_9503), .Z(net_9504) );
CLKBUF_X2 inst_12461 ( .A(net_12159), .Z(net_12309) );
CLKBUF_X2 inst_16390 ( .A(net_16237), .Z(net_16238) );
CLKBUF_X2 inst_9914 ( .A(net_9761), .Z(net_9762) );
CLKBUF_X2 inst_18402 ( .A(net_12249), .Z(net_18250) );
CLKBUF_X2 inst_13205 ( .A(net_13052), .Z(net_13053) );
SDFFR_X2 inst_2203 ( .QN(net_8906), .SE(net_6144), .D(net_2787), .SI(net_2786), .CK(net_17571), .RN(x6501) );
AOI22_X2 inst_8139 ( .B1(net_8186), .A1(net_7676), .B2(net_6099), .A2(net_4399), .ZN(net_4011) );
CLKBUF_X2 inst_13180 ( .A(net_13027), .Z(net_13028) );
CLKBUF_X2 inst_18948 ( .A(net_15411), .Z(net_18796) );
CLKBUF_X2 inst_10495 ( .A(net_10342), .Z(net_10343) );
CLKBUF_X2 inst_14413 ( .A(net_10134), .Z(net_14261) );
CLKBUF_X2 inst_17874 ( .A(net_16720), .Z(net_17722) );
SDFF_X2 inst_1930 ( .SI(net_8058), .Q(net_8058), .D(net_2589), .SE(net_2508), .CK(net_15571) );
CLKBUF_X2 inst_15002 ( .A(net_14849), .Z(net_14850) );
SDFF_X2 inst_577 ( .Q(net_8843), .D(net_8843), .SE(net_3964), .SI(net_3953), .CK(net_10268) );
INV_X4 inst_5536 ( .A(net_1807), .ZN(net_653) );
CLKBUF_X2 inst_12305 ( .A(net_12152), .Z(net_12153) );
CLKBUF_X2 inst_13497 ( .A(net_13344), .Z(net_13345) );
MUX2_X2 inst_4975 ( .A(net_9035), .Z(net_3957), .B(net_3581), .S(net_622) );
CLKBUF_X2 inst_15269 ( .A(net_12155), .Z(net_15117) );
DFF_X1 inst_6760 ( .Q(net_7540), .D(net_4612), .CK(net_11975) );
CLKBUF_X2 inst_17233 ( .A(net_17080), .Z(net_17081) );
NAND3_X2 inst_3938 ( .ZN(net_4936), .A1(net_4688), .A3(net_4681), .A2(net_4484) );
OR2_X2 inst_2865 ( .A2(net_6343), .ZN(net_5940), .A1(net_5714) );
INV_X4 inst_5986 ( .A(net_5977), .ZN(x3561) );
CLKBUF_X2 inst_14933 ( .A(net_14780), .Z(net_14781) );
NAND2_X2 inst_4891 ( .A2(net_7375), .ZN(net_705), .A1(net_164) );
CLKBUF_X2 inst_14520 ( .A(net_14367), .Z(net_14368) );
DFFR_X1 inst_7460 ( .Q(net_7441), .D(net_6189), .CK(net_12854), .RN(x6501) );
CLKBUF_X2 inst_11016 ( .A(net_10167), .Z(net_10864) );
CLKBUF_X2 inst_11092 ( .A(net_9513), .Z(net_10940) );
INV_X2 inst_6264 ( .A(net_8243), .ZN(net_4633) );
CLKBUF_X2 inst_17111 ( .A(net_16958), .Z(net_16959) );
CLKBUF_X2 inst_17384 ( .A(net_17231), .Z(net_17232) );
CLKBUF_X2 inst_14556 ( .A(net_13063), .Z(net_14404) );
DFFR_X2 inst_7040 ( .QN(net_7515), .D(net_4844), .CK(net_13604), .RN(x6501) );
NAND2_X2 inst_4905 ( .A2(net_8267), .A1(net_6149), .ZN(net_611) );
CLKBUF_X2 inst_18350 ( .A(net_18197), .Z(net_18198) );
CLKBUF_X2 inst_17855 ( .A(net_17702), .Z(net_17703) );
XOR2_X2 inst_63 ( .Z(net_928), .A(net_927), .B(net_643) );
AOI22_X2 inst_7968 ( .B1(net_8093), .A1(net_7753), .B2(net_6108), .A2(net_6096), .ZN(net_4161) );
SDFF_X2 inst_1233 ( .Q(net_7830), .D(net_7830), .SE(net_2730), .SI(net_2717), .CK(net_14197) );
INV_X4 inst_5469 ( .A(net_1028), .ZN(net_829) );
OAI22_X2 inst_2924 ( .A2(net_4922), .B1(net_3162), .ZN(net_2938), .B2(net_2888), .A1(net_1882) );
CLKBUF_X2 inst_10445 ( .A(net_10292), .Z(net_10293) );
CLKBUF_X2 inst_11117 ( .A(net_10964), .Z(net_10965) );
SDFF_X2 inst_2006 ( .SI(net_7801), .Q(net_7801), .D(net_2660), .SE(net_2459), .CK(net_16964) );
CLKBUF_X2 inst_10337 ( .A(net_10184), .Z(net_10185) );
SDFFR_X2 inst_2619 ( .Q(net_7376), .D(net_7376), .SE(net_1136), .CK(net_18623), .RN(x6501), .SI(x4771) );
CLKBUF_X2 inst_15625 ( .A(net_11888), .Z(net_15473) );
DFFR_X2 inst_7057 ( .QN(net_7487), .D(net_4773), .CK(net_16669), .RN(x6501) );
SDFF_X2 inst_2033 ( .SI(net_7795), .Q(net_7795), .D(net_2749), .SE(net_2459), .CK(net_14237) );
NOR2_X2 inst_3465 ( .A1(net_3023), .ZN(net_2488), .A2(net_2303) );
CLKBUF_X2 inst_14131 ( .A(net_9238), .Z(net_13979) );
AOI22_X2 inst_7850 ( .A2(net_5595), .ZN(net_4657), .B2(net_4388), .B1(net_2626), .A1(net_320) );
SDFFR_X2 inst_2559 ( .Q(net_6385), .D(net_6385), .SE(net_2147), .SI(net_2129), .CK(net_18239), .RN(x6501) );
CLKBUF_X2 inst_13336 ( .A(net_13183), .Z(net_13184) );
CLKBUF_X2 inst_13898 ( .A(net_13745), .Z(net_13746) );
CLKBUF_X2 inst_16551 ( .A(net_16398), .Z(net_16399) );
CLKBUF_X2 inst_12039 ( .A(net_11886), .Z(net_11887) );
CLKBUF_X2 inst_10201 ( .A(net_10048), .Z(net_10049) );
DFFR_X2 inst_6997 ( .QN(net_6308), .D(net_5850), .CK(net_14224), .RN(x6501) );
AOI22_X2 inst_8386 ( .B1(net_8561), .A1(net_8450), .A2(net_6263), .B2(net_6262), .ZN(net_3662) );
AOI221_X2 inst_8837 ( .C1(net_8174), .B1(net_7732), .C2(net_6101), .B2(net_6095), .ZN(net_6023), .A(net_4290) );
INV_X4 inst_6125 ( .A(net_6374), .ZN(net_683) );
SDFF_X2 inst_1269 ( .Q(net_8102), .D(net_8102), .SI(net_2717), .SE(net_2707), .CK(net_13792) );
CLKBUF_X2 inst_12657 ( .A(net_12504), .Z(net_12505) );
CLKBUF_X2 inst_13575 ( .A(net_13422), .Z(net_13423) );
CLKBUF_X2 inst_14768 ( .A(net_14615), .Z(net_14616) );
CLKBUF_X2 inst_18653 ( .A(net_11955), .Z(net_18501) );
DFFR_X2 inst_7202 ( .D(net_2356), .QN(net_227), .CK(net_17795), .RN(x6501) );
CLKBUF_X2 inst_18301 ( .A(net_18148), .Z(net_18149) );
NOR4_X2 inst_3241 ( .ZN(net_1647), .A1(net_1245), .A3(net_1239), .A2(net_1042), .A4(net_1019) );
CLKBUF_X2 inst_17253 ( .A(net_17100), .Z(net_17101) );
CLKBUF_X2 inst_11842 ( .A(net_11689), .Z(net_11690) );
SDFF_X2 inst_1620 ( .Q(net_8163), .D(net_8163), .SI(net_2719), .SE(net_2538), .CK(net_18786) );
MUX2_X2 inst_4958 ( .A(net_7376), .S(net_2376), .Z(net_2365), .B(net_900) );
CLKBUF_X2 inst_16376 ( .A(net_16223), .Z(net_16224) );
CLKBUF_X2 inst_13344 ( .A(net_11978), .Z(net_13192) );
CLKBUF_X2 inst_10572 ( .A(net_10419), .Z(net_10420) );
SDFF_X2 inst_347 ( .SI(net_8470), .Q(net_8470), .SE(net_3983), .D(net_3954), .CK(net_10087) );
INV_X4 inst_5438 ( .ZN(net_823), .A(net_822) );
CLKBUF_X2 inst_11600 ( .A(net_10267), .Z(net_11448) );
SDFF_X2 inst_755 ( .Q(net_8796), .D(net_8796), .SI(net_3958), .SE(net_3879), .CK(net_13172) );
SDFF_X2 inst_1724 ( .SI(net_7280), .Q(net_7057), .D(net_7057), .SE(net_6280), .CK(net_19024) );
AOI22_X2 inst_7918 ( .A1(net_8994), .A2(net_5456), .B2(net_5260), .ZN(net_4464), .B1(net_3203) );
INV_X4 inst_5855 ( .A(net_7581), .ZN(net_755) );
NAND2_X2 inst_4505 ( .A2(net_6272), .ZN(net_4361), .A1(net_4360) );
CLKBUF_X2 inst_13149 ( .A(net_9248), .Z(net_12997) );
SDFFR_X2 inst_2610 ( .Q(net_7382), .D(net_7382), .SE(net_1136), .CK(net_18651), .RN(x6501), .SI(x4701) );
AOI221_X2 inst_8819 ( .C1(net_7178), .B2(net_6429), .C2(net_5655), .B1(net_5654), .A(net_4905), .ZN(net_4679) );
SDFF_X2 inst_1043 ( .SI(net_7335), .Q(net_6709), .D(net_6709), .SE(net_3125), .CK(net_9760) );
NAND2_X4 inst_4030 ( .A1(net_6200), .ZN(net_6087), .A2(net_2657) );
CLKBUF_X2 inst_12327 ( .A(net_10589), .Z(net_12175) );
DFFR_X2 inst_7230 ( .QN(net_7359), .D(net_2275), .CK(net_11823), .RN(x6501) );
CLKBUF_X2 inst_9234 ( .A(net_9081), .Z(net_9082) );
SDFF_X2 inst_1792 ( .D(net_7273), .SI(net_6890), .Q(net_6890), .SE(net_6284), .CK(net_17379) );
CLKBUF_X2 inst_9769 ( .A(net_9552), .Z(net_9617) );
NAND2_X2 inst_4426 ( .A1(net_6864), .A2(net_5016), .ZN(net_5001) );
INV_X4 inst_6017 ( .A(net_7400), .ZN(net_716) );
CLKBUF_X2 inst_10231 ( .A(net_10078), .Z(net_10079) );
NOR2_X2 inst_3353 ( .ZN(net_5572), .A1(net_5416), .A2(net_5415) );
NAND4_X2 inst_3634 ( .ZN(net_5331), .A2(net_4969), .A1(net_4806), .A4(net_4771), .A3(net_4576) );
CLKBUF_X2 inst_12877 ( .A(net_12724), .Z(net_12725) );
NAND2_X2 inst_4598 ( .ZN(net_2947), .A2(net_2773), .A1(net_1276) );
NAND2_X2 inst_4681 ( .ZN(net_2317), .A1(net_2070), .A2(net_2069) );
CLKBUF_X2 inst_9772 ( .A(net_9080), .Z(net_9620) );
CLKBUF_X2 inst_11204 ( .A(net_10657), .Z(net_11052) );
CLKBUF_X2 inst_16157 ( .A(net_13616), .Z(net_16005) );
CLKBUF_X2 inst_18805 ( .A(net_18652), .Z(net_18653) );
CLKBUF_X2 inst_18490 ( .A(net_18337), .Z(net_18338) );
OAI21_X2 inst_3145 ( .A(net_2304), .ZN(net_2030), .B2(net_1935), .B1(net_1751) );
INV_X4 inst_5144 ( .ZN(net_3358), .A(net_3301) );
SDFF_X2 inst_648 ( .Q(net_8419), .D(net_8419), .SI(net_3962), .SE(net_3934), .CK(net_10153) );
CLKBUF_X2 inst_10600 ( .A(net_10447), .Z(net_10448) );
AOI22_X2 inst_7857 ( .A2(net_5595), .B2(net_4881), .ZN(net_4650), .A1(net_327), .B1(net_245) );
CLKBUF_X2 inst_13718 ( .A(net_13565), .Z(net_13566) );
CLKBUF_X2 inst_16363 ( .A(net_16210), .Z(net_16211) );
XNOR2_X2 inst_270 ( .B(net_1121), .ZN(net_1050), .A(net_548) );
SDFF_X2 inst_1901 ( .D(net_7294), .SI(net_7031), .Q(net_7031), .SE(net_6277), .CK(net_17662) );
NAND2_X2 inst_4104 ( .ZN(net_5428), .A1(net_5152), .A2(net_5151) );
CLKBUF_X2 inst_11826 ( .A(net_11673), .Z(net_11674) );
AOI222_X1 inst_8608 ( .B2(net_6756), .C2(net_6198), .B1(net_5835), .ZN(net_5815), .A2(net_3114), .A1(net_837), .C1(x3604) );
SDFFR_X2 inst_2552 ( .QN(net_6358), .SE(net_2147), .D(net_2132), .SI(net_1866), .CK(net_17402), .RN(x6501) );
CLKBUF_X2 inst_18914 ( .A(net_18761), .Z(net_18762) );
SDFF_X2 inst_631 ( .SI(net_8544), .Q(net_8544), .SE(net_3979), .D(net_3954), .CK(net_10063) );
CLKBUF_X2 inst_11809 ( .A(net_11656), .Z(net_11657) );
CLKBUF_X2 inst_18712 ( .A(net_18559), .Z(net_18560) );
INV_X2 inst_6427 ( .A(net_841), .ZN(net_735) );
CLKBUF_X2 inst_15070 ( .A(net_13019), .Z(net_14918) );
NAND4_X2 inst_3674 ( .A4(net_6059), .A1(net_6058), .ZN(net_4591), .A2(net_4048), .A3(net_4047) );
CLKBUF_X2 inst_12835 ( .A(net_12682), .Z(net_12683) );
CLKBUF_X2 inst_11346 ( .A(net_11193), .Z(net_11194) );
CLKBUF_X2 inst_13505 ( .A(net_13352), .Z(net_13353) );
CLKBUF_X2 inst_13789 ( .A(net_13636), .Z(net_13637) );
NAND3_X2 inst_3995 ( .A3(net_4320), .ZN(net_1732), .A2(net_1522), .A1(net_1372) );
INV_X4 inst_5074 ( .ZN(net_5854), .A(net_5806) );
CLKBUF_X2 inst_19198 ( .A(net_19045), .Z(net_19046) );
XOR2_X1 inst_102 ( .A(net_7649), .B(net_3082), .Z(net_1182) );
CLKBUF_X2 inst_14749 ( .A(net_13691), .Z(net_14597) );
SDFFR_X2 inst_2527 ( .D(net_7367), .SE(net_2387), .SI(net_282), .Q(net_282), .CK(net_16383), .RN(x6501) );
NOR3_X2 inst_3277 ( .ZN(net_2814), .A1(net_2400), .A3(net_2398), .A2(net_1461) );
CLKBUF_X2 inst_12042 ( .A(net_11889), .Z(net_11890) );
SDFFR_X1 inst_2786 ( .D(net_7376), .Q(net_7273), .SI(net_1866), .SE(net_1327), .CK(net_17409), .RN(x6501) );
INV_X4 inst_5352 ( .A(net_1921), .ZN(net_1177) );
SDFF_X2 inst_1224 ( .Q(net_7943), .D(net_7943), .SE(net_2755), .SI(net_2585), .CK(net_18590) );
CLKBUF_X2 inst_10043 ( .A(net_9511), .Z(net_9891) );
CLKBUF_X2 inst_11045 ( .A(net_10892), .Z(net_10893) );
CLKBUF_X2 inst_16040 ( .A(net_15887), .Z(net_15888) );
NAND3_X2 inst_3905 ( .ZN(net_5633), .A1(net_5562), .A3(net_5496), .A2(net_5374) );
SDFF_X2 inst_1170 ( .D(net_7337), .SI(net_6513), .Q(net_6513), .SE(net_3071), .CK(net_9443) );
AOI21_X2 inst_8929 ( .B2(net_5843), .ZN(net_5682), .A(net_5668), .B1(x378) );
CLKBUF_X2 inst_11797 ( .A(net_10666), .Z(net_11645) );
CLKBUF_X2 inst_16886 ( .A(net_12855), .Z(net_16734) );
CLKBUF_X2 inst_14246 ( .A(net_9180), .Z(net_14094) );
CLKBUF_X2 inst_15219 ( .A(net_15066), .Z(net_15067) );
CLKBUF_X2 inst_11659 ( .A(net_10936), .Z(net_11507) );
AOI221_X2 inst_8752 ( .C2(net_6454), .C1(net_5654), .B2(net_5595), .ZN(net_5594), .A(net_5331), .B1(net_336) );
CLKBUF_X2 inst_17373 ( .A(net_17220), .Z(net_17221) );
SDFF_X2 inst_785 ( .SI(net_8354), .Q(net_8354), .D(net_3957), .SE(net_3880), .CK(net_13237) );
SDFFR_X2 inst_2362 ( .SE(net_2260), .Q(net_368), .D(net_368), .CK(net_11457), .RN(x6501), .SI(x1721) );
CLKBUF_X2 inst_18389 ( .A(net_18236), .Z(net_18237) );
OR2_X4 inst_2856 ( .A1(net_6807), .A2(net_6804), .ZN(net_774) );
CLKBUF_X2 inst_9280 ( .A(net_9127), .Z(net_9128) );
CLKBUF_X2 inst_10417 ( .A(net_10264), .Z(net_10265) );
AOI22_X2 inst_7945 ( .B1(net_8158), .A1(net_7716), .B2(net_6101), .A2(net_6095), .ZN(net_6000) );
SDFF_X2 inst_527 ( .Q(net_8883), .D(net_8883), .SI(net_3951), .SE(net_3936), .CK(net_10604) );
XNOR2_X2 inst_226 ( .ZN(net_1362), .B(net_1361), .A(net_531) );
SDFF_X2 inst_1180 ( .SI(net_7334), .Q(net_6609), .D(net_6609), .SE(net_3069), .CK(net_9742) );
INV_X4 inst_5509 ( .ZN(net_860), .A(net_689) );
CLKBUF_X2 inst_19066 ( .A(net_18913), .Z(net_18914) );
AOI22_X2 inst_8223 ( .B1(net_8685), .A1(net_8648), .ZN(net_6248), .B2(net_6109), .A2(net_3857) );
CLKBUF_X2 inst_13861 ( .A(net_13708), .Z(net_13709) );
CLKBUF_X2 inst_11232 ( .A(net_11079), .Z(net_11080) );
XNOR2_X2 inst_212 ( .ZN(net_1449), .B(net_1308), .A(net_1307) );
CLKBUF_X2 inst_11688 ( .A(net_9246), .Z(net_11536) );
SDFFR_X1 inst_2732 ( .SI(net_9045), .Q(net_9045), .D(net_7474), .SE(net_3208), .CK(net_12212), .RN(x6501) );
CLKBUF_X2 inst_16682 ( .A(net_16529), .Z(net_16530) );
INV_X2 inst_6321 ( .ZN(net_3342), .A(net_3287) );
CLKBUF_X2 inst_9323 ( .A(net_9170), .Z(net_9171) );
CLKBUF_X2 inst_15293 ( .A(net_15140), .Z(net_15141) );
CLKBUF_X2 inst_18627 ( .A(net_9702), .Z(net_18475) );
CLKBUF_X2 inst_18771 ( .A(net_18618), .Z(net_18619) );
CLKBUF_X2 inst_10013 ( .A(net_9804), .Z(net_9861) );
INV_X4 inst_5431 ( .A(net_7401), .ZN(net_1149) );
AOI22_X2 inst_8330 ( .B1(net_8587), .A1(net_8476), .A2(net_6263), .B2(net_6262), .ZN(net_3716) );
CLKBUF_X2 inst_14638 ( .A(net_9873), .Z(net_14486) );
OAI221_X2 inst_2966 ( .ZN(net_2654), .B2(net_2650), .C2(net_2649), .A(net_2481), .B1(net_1844), .C1(net_1043) );
NOR4_X2 inst_3246 ( .ZN(net_1556), .A1(net_1050), .A2(net_1008), .A4(net_984), .A3(net_819) );
NAND2_X2 inst_4904 ( .A2(net_7395), .ZN(net_615), .A1(net_184) );
CLKBUF_X2 inst_16440 ( .A(net_16287), .Z(net_16288) );
CLKBUF_X2 inst_19059 ( .A(net_18906), .Z(net_18907) );
CLKBUF_X2 inst_16803 ( .A(net_16650), .Z(net_16651) );
NAND2_X2 inst_4887 ( .A2(net_7163), .A1(net_7162), .ZN(net_710) );
CLKBUF_X2 inst_11272 ( .A(net_11119), .Z(net_11120) );
SDFFR_X2 inst_2381 ( .SE(net_2260), .Q(net_336), .D(net_336), .CK(net_9291), .RN(x6501), .SI(x2355) );
INV_X4 inst_5823 ( .A(net_6398), .ZN(net_2832) );
CLKBUF_X2 inst_11538 ( .A(net_9766), .Z(net_11386) );
CLKBUF_X2 inst_16059 ( .A(net_13980), .Z(net_15907) );
CLKBUF_X2 inst_11284 ( .A(net_11131), .Z(net_11132) );
CLKBUF_X2 inst_16922 ( .A(net_15105), .Z(net_16770) );
CLKBUF_X2 inst_18947 ( .A(net_18794), .Z(net_18795) );
SDFF_X2 inst_454 ( .SI(net_8456), .Q(net_8456), .SE(net_3983), .D(net_3962), .CK(net_10191) );
CLKBUF_X2 inst_13753 ( .A(net_13600), .Z(net_13601) );
CLKBUF_X2 inst_13947 ( .A(net_13794), .Z(net_13795) );
CLKBUF_X2 inst_14299 ( .A(net_12276), .Z(net_14147) );
CLKBUF_X2 inst_18719 ( .A(net_18566), .Z(net_18567) );
AOI22_X2 inst_8251 ( .B1(net_8688), .A1(net_8651), .B2(net_6109), .A2(net_3857), .ZN(net_3785) );
CLKBUF_X2 inst_15475 ( .A(net_13150), .Z(net_15323) );
CLKBUF_X2 inst_17035 ( .A(net_16674), .Z(net_16883) );
AOI22_X2 inst_7899 ( .A2(net_4553), .ZN(net_4530), .B1(net_2931), .B2(net_1634), .A1(net_1606) );
CLKBUF_X2 inst_16175 ( .A(net_16022), .Z(net_16023) );
CLKBUF_X2 inst_11130 ( .A(net_9348), .Z(net_10978) );
CLKBUF_X2 inst_11067 ( .A(net_9442), .Z(net_10915) );
DFFR_X2 inst_6990 ( .QN(net_5970), .D(net_5890), .CK(net_11552), .RN(x6501) );
CLKBUF_X2 inst_13622 ( .A(net_13469), .Z(net_13470) );
CLKBUF_X2 inst_12974 ( .A(net_10015), .Z(net_12822) );
SDFFR_X2 inst_2419 ( .D(net_2684), .SE(net_2683), .SI(net_466), .Q(net_466), .CK(net_16909), .RN(x6501) );
CLKBUF_X2 inst_14793 ( .A(net_14640), .Z(net_14641) );
CLKBUF_X2 inst_9484 ( .A(net_9211), .Z(net_9332) );
CLKBUF_X2 inst_11612 ( .A(net_9433), .Z(net_11460) );
CLKBUF_X2 inst_17996 ( .A(net_17843), .Z(net_17844) );
INV_X8 inst_5041 ( .ZN(net_6101), .A(net_3577) );
SDFF_X2 inst_1428 ( .SI(net_7288), .Q(net_7065), .D(net_7065), .SE(net_6280), .CK(net_17714) );
CLKBUF_X2 inst_11089 ( .A(net_10936), .Z(net_10937) );
CLKBUF_X2 inst_16467 ( .A(net_15196), .Z(net_16315) );
CLKBUF_X2 inst_9456 ( .A(net_9303), .Z(net_9304) );
SDFFR_X1 inst_2739 ( .SI(net_9021), .Q(net_9021), .D(net_7450), .SE(net_3208), .CK(net_10099), .RN(x6501) );
CLKBUF_X2 inst_12691 ( .A(net_11707), .Z(net_12539) );
SDFF_X2 inst_1046 ( .SI(net_7324), .Q(net_6698), .D(net_6698), .SE(net_3125), .CK(net_9860) );
INV_X4 inst_5955 ( .A(net_8957), .ZN(net_1757) );
NAND2_X2 inst_4355 ( .A1(net_7069), .A2(net_5162), .ZN(net_5102) );
CLKBUF_X2 inst_10152 ( .A(net_9999), .Z(net_10000) );
INV_X4 inst_5426 ( .A(net_7399), .ZN(net_1129) );
INV_X2 inst_6206 ( .ZN(net_5504), .A(net_5405) );
CLKBUF_X2 inst_9515 ( .A(net_9362), .Z(net_9363) );
CLKBUF_X2 inst_16859 ( .A(net_11774), .Z(net_16707) );
CLKBUF_X2 inst_16454 ( .A(net_16301), .Z(net_16302) );
SDFF_X2 inst_909 ( .SI(net_8727), .Q(net_8727), .SE(net_6195), .D(net_3942), .CK(net_12574) );
CLKBUF_X2 inst_17393 ( .A(net_17240), .Z(net_17241) );
SDFFR_X2 inst_2484 ( .Q(net_8984), .D(net_8984), .SI(net_2614), .SE(net_2562), .CK(net_13921), .RN(x6501) );
INV_X4 inst_5758 ( .A(net_7579), .ZN(net_626) );
CLKBUF_X2 inst_9927 ( .A(net_9225), .Z(net_9775) );
CLKBUF_X2 inst_19148 ( .A(net_18995), .Z(net_18996) );
INV_X2 inst_6494 ( .A(net_6352), .ZN(net_2128) );
OAI22_X2 inst_2919 ( .ZN(net_3257), .A2(net_3147), .B2(net_3146), .A1(net_1693), .B1(net_604) );
SDFF_X2 inst_1872 ( .D(net_7275), .SI(net_6972), .Q(net_6972), .SE(net_6283), .CK(net_14618) );
INV_X8 inst_5039 ( .ZN(net_6096), .A(net_3530) );
CLKBUF_X2 inst_10795 ( .A(net_10642), .Z(net_10643) );
CLKBUF_X2 inst_10827 ( .A(net_10674), .Z(net_10675) );
CLKBUF_X2 inst_12003 ( .A(net_11850), .Z(net_11851) );
CLKBUF_X2 inst_15917 ( .A(net_15764), .Z(net_15765) );
NAND2_X4 inst_4028 ( .ZN(net_3123), .A2(net_2940), .A1(net_2905) );
AOI22_X2 inst_8478 ( .B1(net_6675), .A1(net_6642), .A2(net_6213), .B2(net_6138), .ZN(net_3462) );
CLKBUF_X2 inst_16658 ( .A(net_16505), .Z(net_16506) );
CLKBUF_X2 inst_17640 ( .A(net_17487), .Z(net_17488) );
CLKBUF_X2 inst_17608 ( .A(net_11352), .Z(net_17456) );
CLKBUF_X2 inst_17136 ( .A(net_16983), .Z(net_16984) );
CLKBUF_X2 inst_16083 ( .A(net_15930), .Z(net_15931) );
CLKBUF_X2 inst_13556 ( .A(net_13403), .Z(net_13404) );
CLKBUF_X2 inst_18200 ( .A(net_18047), .Z(net_18048) );
OAI21_X2 inst_3119 ( .ZN(net_2305), .A(net_2304), .B2(net_2241), .B1(net_2124) );
NAND4_X2 inst_3777 ( .ZN(net_4244), .A1(net_3724), .A2(net_3723), .A3(net_3722), .A4(net_3721) );
INV_X4 inst_5138 ( .ZN(net_3570), .A(net_3563) );
CLKBUF_X2 inst_18109 ( .A(net_11738), .Z(net_17957) );
XOR2_X2 inst_29 ( .A(net_7585), .B(net_3227), .Z(net_1223) );
CLKBUF_X2 inst_14515 ( .A(net_14362), .Z(net_14363) );
CLKBUF_X2 inst_9900 ( .A(net_9656), .Z(net_9748) );
DFFS_X1 inst_6937 ( .D(net_6145), .CK(net_13653), .SN(x6501), .Q(x719) );
AOI22_X2 inst_8469 ( .B1(net_6739), .A1(net_6706), .B2(net_6202), .A2(net_3520), .ZN(net_3471) );
AOI22_X2 inst_7782 ( .A1(net_5268), .ZN(net_4869), .A2(net_4633), .B2(net_4388), .B1(net_2632) );
CLKBUF_X2 inst_9713 ( .A(net_9397), .Z(net_9561) );
CLKBUF_X2 inst_16471 ( .A(net_16318), .Z(net_16319) );
SDFFR_X2 inst_2152 ( .Q(net_8277), .D(net_8277), .SI(net_8273), .SE(net_2996), .CK(net_18446), .RN(x6501) );
NAND3_X2 inst_3947 ( .A3(net_6211), .ZN(net_4325), .A1(net_4324), .A2(net_1129) );
CLKBUF_X2 inst_10540 ( .A(net_10387), .Z(net_10388) );
CLKBUF_X2 inst_16232 ( .A(net_14150), .Z(net_16080) );
AOI22_X2 inst_7740 ( .B1(net_6960), .A1(net_6920), .ZN(net_5448), .A2(net_5443), .B2(net_5442) );
CLKBUF_X2 inst_13270 ( .A(net_12775), .Z(net_13118) );
CLKBUF_X2 inst_15712 ( .A(net_15247), .Z(net_15560) );
CLKBUF_X2 inst_10590 ( .A(net_10437), .Z(net_10438) );
CLKBUF_X2 inst_11152 ( .A(net_10999), .Z(net_11000) );
CLKBUF_X2 inst_12775 ( .A(net_12622), .Z(net_12623) );
INV_X2 inst_6207 ( .ZN(net_5503), .A(net_5401) );
CLKBUF_X2 inst_11396 ( .A(net_11243), .Z(net_11244) );
SDFF_X2 inst_538 ( .Q(net_8679), .D(net_8679), .SI(net_3945), .SE(net_3935), .CK(net_11092) );
AOI22_X2 inst_8344 ( .B1(net_8589), .A1(net_8478), .A2(net_6263), .B2(net_6262), .ZN(net_3703) );
CLKBUF_X2 inst_16277 ( .A(net_16124), .Z(net_16125) );
NAND2_X2 inst_4537 ( .A2(net_3373), .ZN(net_3372), .A1(net_3371) );
INV_X4 inst_5280 ( .A(net_2318), .ZN(net_1885) );
XOR2_X2 inst_35 ( .B(net_2758), .A(net_2667), .Z(net_1185) );
NAND2_X2 inst_4765 ( .A2(net_6169), .A1(net_2520), .ZN(net_1693) );
AOI21_X2 inst_8890 ( .B2(net_5871), .ZN(net_5806), .A(net_5805), .B1(net_2689) );
CLKBUF_X2 inst_10599 ( .A(net_10446), .Z(net_10447) );
CLKBUF_X2 inst_11146 ( .A(net_9714), .Z(net_10994) );
SDFFR_X2 inst_2600 ( .D(net_7373), .Q(net_7270), .SI(net_1856), .SE(net_1327), .CK(net_14684), .RN(x6501) );
CLKBUF_X2 inst_14158 ( .A(net_14005), .Z(net_14006) );
CLKBUF_X2 inst_16990 ( .A(net_12206), .Z(net_16838) );
SDFFR_X2 inst_2274 ( .SI(net_7385), .SE(net_2814), .Q(net_244), .D(net_244), .CK(net_17540), .RN(x6501) );
INV_X4 inst_5178 ( .ZN(net_2941), .A(net_2911) );
CLKBUF_X2 inst_10055 ( .A(net_9902), .Z(net_9903) );
CLKBUF_X2 inst_16671 ( .A(net_16518), .Z(net_16519) );
SDFF_X2 inst_695 ( .Q(net_8868), .D(net_8868), .SI(net_3944), .SE(net_3936), .CK(net_12264) );
CLKBUF_X2 inst_19016 ( .A(net_18863), .Z(net_18864) );
NAND2_X4 inst_4038 ( .ZN(net_6089), .A1(net_2403), .A2(net_2324) );
INV_X4 inst_5492 ( .A(net_1806), .ZN(net_721) );
CLKBUF_X2 inst_10606 ( .A(net_9440), .Z(net_10454) );
CLKBUF_X2 inst_10663 ( .A(net_10510), .Z(net_10511) );
CLKBUF_X2 inst_14001 ( .A(net_13848), .Z(net_13849) );
DFFS_X2 inst_6877 ( .QN(net_6458), .D(net_3347), .CK(net_17926), .SN(x6501) );
CLKBUF_X2 inst_10782 ( .A(net_10629), .Z(net_10630) );
CLKBUF_X2 inst_14376 ( .A(net_14223), .Z(net_14224) );
INV_X4 inst_6154 ( .A(net_6183), .ZN(net_6182) );
NOR2_X2 inst_3559 ( .ZN(net_3308), .A2(net_1342), .A1(net_496) );
CLKBUF_X2 inst_17790 ( .A(net_14995), .Z(net_17638) );
CLKBUF_X2 inst_17306 ( .A(net_17153), .Z(net_17154) );
INV_X4 inst_5720 ( .A(net_7252), .ZN(net_1951) );
CLKBUF_X2 inst_12277 ( .A(net_12124), .Z(net_12125) );
CLKBUF_X2 inst_17688 ( .A(net_17535), .Z(net_17536) );
CLKBUF_X2 inst_9449 ( .A(net_9296), .Z(net_9297) );
CLKBUF_X2 inst_17386 ( .A(net_17233), .Z(net_17234) );
DFFR_X2 inst_7183 ( .QN(net_5954), .D(net_2485), .CK(net_16295), .RN(x6501) );
AOI22_X2 inst_8328 ( .B1(net_8772), .A1(net_8402), .A2(net_3867), .B2(net_3866), .ZN(net_3718) );
CLKBUF_X2 inst_11772 ( .A(net_11619), .Z(net_11620) );
CLKBUF_X2 inst_12790 ( .A(net_12637), .Z(net_12638) );
CLKBUF_X2 inst_16315 ( .A(net_16162), .Z(net_16163) );
INV_X4 inst_6001 ( .A(net_7403), .ZN(net_664) );
DFFR_X2 inst_7004 ( .D(net_5873), .CK(net_9229), .RN(x6501), .Q(x2355) );
CLKBUF_X2 inst_12506 ( .A(net_12353), .Z(net_12354) );
CLKBUF_X2 inst_18268 ( .A(net_18115), .Z(net_18116) );
CLKBUF_X2 inst_16995 ( .A(net_16842), .Z(net_16843) );
AOI22_X2 inst_8193 ( .B1(net_8828), .A1(net_8347), .A2(net_6265), .B2(net_6253), .ZN(net_6074) );
CLKBUF_X2 inst_19102 ( .A(net_14131), .Z(net_18950) );
CLKBUF_X2 inst_14086 ( .A(net_10583), .Z(net_13934) );
CLKBUF_X2 inst_11646 ( .A(net_10738), .Z(net_11494) );
CLKBUF_X2 inst_10751 ( .A(net_10598), .Z(net_10599) );
CLKBUF_X2 inst_11525 ( .A(net_11372), .Z(net_11373) );
CLKBUF_X2 inst_10666 ( .A(net_9515), .Z(net_10514) );
INV_X2 inst_6592 ( .A(net_6123), .ZN(net_6122) );
DFFR_X2 inst_7209 ( .D(net_2360), .QN(net_220), .CK(net_17474), .RN(x6501) );
CLKBUF_X2 inst_14865 ( .A(net_14712), .Z(net_14713) );
INV_X4 inst_5217 ( .ZN(net_2403), .A(net_2321) );
AOI22_X2 inst_8069 ( .B1(net_8038), .A1(net_8004), .B2(net_6102), .A2(net_6097), .ZN(net_4074) );
CLKBUF_X2 inst_15307 ( .A(net_15154), .Z(net_15155) );
NAND2_X2 inst_4600 ( .A2(net_2897), .ZN(net_2894), .A1(net_2770) );
NAND3_X4 inst_3872 ( .A3(net_7344), .ZN(net_6147), .A1(net_6079), .A2(net_2251) );
DFFS_X1 inst_6923 ( .D(net_6145), .CK(net_13658), .SN(x6501), .Q(x808) );
CLKBUF_X2 inst_9273 ( .A(net_9110), .Z(net_9121) );
CLKBUF_X2 inst_11574 ( .A(net_11421), .Z(net_11422) );
CLKBUF_X2 inst_17067 ( .A(net_11445), .Z(net_16915) );
CLKBUF_X2 inst_10227 ( .A(net_10074), .Z(net_10075) );
CLKBUF_X2 inst_17849 ( .A(net_12144), .Z(net_17697) );
SDFF_X2 inst_1411 ( .SI(net_7284), .Q(net_7101), .D(net_7101), .SE(net_6278), .CK(net_16239) );
XNOR2_X2 inst_149 ( .ZN(net_2108), .B(net_1826), .A(net_1823) );
CLKBUF_X2 inst_11028 ( .A(net_10875), .Z(net_10876) );
CLKBUF_X2 inst_12527 ( .A(net_12374), .Z(net_12375) );
CLKBUF_X2 inst_18048 ( .A(net_17895), .Z(net_17896) );
AOI221_X2 inst_8854 ( .B1(net_8584), .C1(net_8473), .C2(net_6263), .B2(net_6262), .ZN(net_6229), .A(net_4247) );
DFFS_X1 inst_6924 ( .D(net_6145), .CK(net_16376), .SN(x6501), .Q(x815) );
CLKBUF_X2 inst_18134 ( .A(net_16198), .Z(net_17982) );
CLKBUF_X2 inst_9542 ( .A(net_9389), .Z(net_9390) );
AOI22_X2 inst_7771 ( .B1(net_6998), .A1(net_6958), .A2(net_5443), .B2(net_5442), .ZN(net_5319) );
CLKBUF_X2 inst_15608 ( .A(net_15455), .Z(net_15456) );
SDFFR_X2 inst_2320 ( .SE(net_2748), .D(net_2744), .SI(net_461), .Q(net_461), .CK(net_16924), .RN(x6501) );
CLKBUF_X2 inst_15203 ( .A(net_15050), .Z(net_15051) );
CLKBUF_X2 inst_17582 ( .A(net_17429), .Z(net_17430) );
SDFFR_X2 inst_2534 ( .QN(net_6361), .SE(net_2147), .SI(net_1941), .D(net_690), .CK(net_14763), .RN(x6501) );
CLKBUF_X2 inst_17527 ( .A(net_17374), .Z(net_17375) );
INV_X4 inst_5377 ( .A(net_2097), .ZN(net_1377) );
CLKBUF_X2 inst_10775 ( .A(net_10622), .Z(net_10623) );
NAND4_X2 inst_3737 ( .ZN(net_4293), .A1(net_4094), .A2(net_4093), .A3(net_4092), .A4(net_4091) );
SDFF_X2 inst_1636 ( .Q(net_8151), .D(net_8151), .SI(net_2659), .SE(net_2538), .CK(net_18546) );
SDFF_X2 inst_515 ( .Q(net_8869), .D(net_8869), .SI(net_3967), .SE(net_3936), .CK(net_10022) );
AOI22_X2 inst_8501 ( .B1(net_6747), .A1(net_6714), .B2(net_6202), .A2(net_3520), .ZN(net_3439) );
SDFF_X2 inst_1501 ( .SI(net_7859), .Q(net_7859), .D(net_2722), .SE(net_2558), .CK(net_18791) );
DFFR_X2 inst_7278 ( .Q(net_7223), .D(net_2066), .CK(net_15185), .RN(x6501) );
CLKBUF_X2 inst_12242 ( .A(net_9903), .Z(net_12090) );
OAI211_X2 inst_3212 ( .B(net_4685), .A(net_2077), .ZN(net_1999), .C2(net_1998), .C1(net_1692) );
CLKBUF_X2 inst_14982 ( .A(net_12919), .Z(net_14830) );
SDFF_X2 inst_1584 ( .Q(net_8038), .D(net_8038), .SI(net_2715), .SE(net_2545), .CK(net_14172) );
CLKBUF_X2 inst_14183 ( .A(net_14030), .Z(net_14031) );
CLKBUF_X2 inst_9361 ( .A(net_9176), .Z(net_9209) );
AOI22_X2 inst_7933 ( .B1(net_8088), .A1(net_7748), .B2(net_6108), .A2(net_6096), .ZN(net_4192) );
CLKBUF_X2 inst_11023 ( .A(net_10870), .Z(net_10871) );
CLKBUF_X2 inst_15499 ( .A(net_15346), .Z(net_15347) );
AOI22_X2 inst_8129 ( .B1(net_8117), .A1(net_7879), .A2(net_6098), .B2(net_4190), .ZN(net_4020) );
OAI22_X2 inst_2933 ( .B2(net_2299), .A2(net_2187), .ZN(net_2176), .A1(net_2175), .B1(net_1963) );
INV_X2 inst_6467 ( .A(net_7364), .ZN(net_574) );
AOI221_X4 inst_8706 ( .C1(net_8194), .B1(net_7684), .C2(net_6099), .ZN(net_6035), .B2(net_4399), .A(net_4305) );
CLKBUF_X2 inst_14641 ( .A(net_14488), .Z(net_14489) );
SDFFR_X1 inst_2713 ( .D(net_7163), .QN(net_6423), .SE(net_4624), .SI(net_1829), .CK(net_9540), .RN(x6501) );
SDFF_X2 inst_1008 ( .D(net_7320), .SI(net_6628), .Q(net_6628), .SE(net_3123), .CK(net_12112) );
SDFF_X2 inst_559 ( .Q(net_8674), .D(net_8674), .SI(net_3981), .SE(net_3935), .CK(net_12988) );
AOI22_X2 inst_7877 ( .B2(net_4881), .ZN(net_4563), .A2(net_4562), .A1(net_1657), .B1(net_256) );
AOI21_X2 inst_8872 ( .B2(net_6254), .ZN(net_5935), .A(net_5934), .B1(x1039) );
DFF_X1 inst_6725 ( .Q(net_6771), .D(net_5644), .CK(net_9259) );
CLKBUF_X2 inst_9476 ( .A(net_9323), .Z(net_9324) );
CLKBUF_X2 inst_11596 ( .A(net_11354), .Z(net_11444) );
CLKBUF_X2 inst_19012 ( .A(net_10950), .Z(net_18860) );
CLKBUF_X2 inst_9250 ( .A(net_9097), .Z(net_9098) );
CLKBUF_X2 inst_14940 ( .A(net_14787), .Z(net_14788) );
CLKBUF_X2 inst_18933 ( .A(net_18780), .Z(net_18781) );
CLKBUF_X2 inst_16818 ( .A(net_13271), .Z(net_16666) );
NOR2_X2 inst_3405 ( .A2(net_6145), .ZN(net_3876), .A1(net_3322) );
NAND3_X2 inst_3888 ( .ZN(net_5650), .A1(net_5579), .A3(net_5513), .A2(net_5444) );
AOI21_X2 inst_8979 ( .B1(net_7165), .B2(net_2146), .ZN(net_2100), .A(net_2099) );
CLKBUF_X2 inst_12831 ( .A(net_12200), .Z(net_12679) );
CLKBUF_X2 inst_9797 ( .A(net_9644), .Z(net_9645) );
DFFR_X2 inst_7366 ( .Q(net_7336), .CK(net_11703), .D(x12955), .RN(x6501) );
CLKBUF_X2 inst_12221 ( .A(net_12068), .Z(net_12069) );
CLKBUF_X2 inst_15275 ( .A(net_11161), .Z(net_15123) );
NAND2_X2 inst_4334 ( .A1(net_7062), .A2(net_5162), .ZN(net_5123) );
AOI22_X2 inst_8017 ( .A1(net_7963), .B1(net_7793), .A2(net_6092), .B2(net_6091), .ZN(net_4119) );
SDFF_X2 inst_1075 ( .D(net_7324), .SI(net_6500), .Q(net_6500), .SE(net_3071), .CK(net_11322) );
CLKBUF_X2 inst_19038 ( .A(net_18565), .Z(net_18886) );
CLKBUF_X2 inst_9230 ( .A(net_9063), .Z(net_9078) );
CLKBUF_X2 inst_12701 ( .A(net_9414), .Z(net_12549) );
SDFFR_X2 inst_2257 ( .D(net_7388), .SE(net_2797), .SI(net_197), .Q(net_197), .CK(net_17547), .RN(x6501) );
CLKBUF_X2 inst_11504 ( .A(net_10551), .Z(net_11352) );
CLKBUF_X2 inst_11781 ( .A(net_11628), .Z(net_11629) );
CLKBUF_X2 inst_16183 ( .A(net_9173), .Z(net_16031) );
CLKBUF_X2 inst_15278 ( .A(net_10263), .Z(net_15126) );
CLKBUF_X2 inst_13641 ( .A(net_12165), .Z(net_13489) );
CLKBUF_X2 inst_14306 ( .A(net_12441), .Z(net_14154) );
CLKBUF_X2 inst_15553 ( .A(net_15133), .Z(net_15401) );
CLKBUF_X2 inst_15210 ( .A(net_15057), .Z(net_15058) );
INV_X2 inst_6536 ( .A(net_7348), .ZN(net_686) );
INV_X4 inst_6110 ( .A(net_6797), .ZN(net_4373) );
INV_X2 inst_6434 ( .ZN(net_687), .A(net_686) );
SDFF_X2 inst_494 ( .SI(net_8619), .Q(net_8619), .SE(net_3984), .D(net_3975), .CK(net_12546) );
XNOR2_X2 inst_329 ( .B(net_7591), .A(net_7442), .ZN(net_840) );
CLKBUF_X2 inst_17823 ( .A(net_17670), .Z(net_17671) );
INV_X4 inst_5942 ( .A(net_7240), .ZN(net_1943) );
SDFFR_X2 inst_2347 ( .SE(net_2260), .Q(net_316), .D(net_316), .CK(net_10439), .RN(x6501), .SI(x3288) );
CLKBUF_X2 inst_13845 ( .A(net_13692), .Z(net_13693) );
CLKBUF_X2 inst_13085 ( .A(net_12734), .Z(net_12933) );
CLKBUF_X2 inst_17117 ( .A(net_9144), .Z(net_16965) );
CLKBUF_X2 inst_14167 ( .A(net_10913), .Z(net_14015) );
OR2_X2 inst_2894 ( .A2(net_2902), .A1(net_2901), .ZN(net_2770) );
INV_X4 inst_5949 ( .A(net_7413), .ZN(net_1468) );
DFFR_X2 inst_7045 ( .QN(net_8899), .D(net_4895), .CK(net_17640), .RN(x6501) );
INV_X4 inst_6085 ( .ZN(net_2731), .A(net_144) );
CLKBUF_X2 inst_10192 ( .A(net_10039), .Z(net_10040) );
OAI221_X2 inst_2959 ( .C2(net_8248), .B1(net_7591), .B2(net_4971), .C1(net_4928), .ZN(net_4844), .A(net_3333) );
CLKBUF_X2 inst_15130 ( .A(net_14977), .Z(net_14978) );
CLKBUF_X2 inst_18474 ( .A(net_16981), .Z(net_18322) );
CLKBUF_X2 inst_13906 ( .A(net_13753), .Z(net_13754) );
CLKBUF_X2 inst_19194 ( .A(net_18448), .Z(net_19042) );
SDFF_X2 inst_1683 ( .SI(net_7283), .Q(net_7060), .D(net_7060), .SE(net_6280), .CK(net_16211) );
CLKBUF_X2 inst_10714 ( .A(net_10561), .Z(net_10562) );
NAND3_X4 inst_3865 ( .A3(net_6259), .A2(net_6194), .ZN(net_4902), .A1(net_4901) );
CLKBUF_X2 inst_18003 ( .A(net_9104), .Z(net_17851) );
CLKBUF_X2 inst_16983 ( .A(net_16830), .Z(net_16831) );
CLKBUF_X2 inst_10459 ( .A(net_9973), .Z(net_10307) );
CLKBUF_X2 inst_13109 ( .A(net_12100), .Z(net_12957) );
CLKBUF_X2 inst_9896 ( .A(net_9743), .Z(net_9744) );
CLKBUF_X2 inst_15099 ( .A(net_14946), .Z(net_14947) );
NOR2_X2 inst_3543 ( .ZN(net_1470), .A2(net_1469), .A1(net_1070) );
CLKBUF_X2 inst_15486 ( .A(net_11080), .Z(net_15334) );
HA_X1 inst_6712 ( .A(net_6460), .B(net_3292), .S(net_1233), .CO(net_1232) );
CLKBUF_X2 inst_10737 ( .A(net_9889), .Z(net_10585) );
CLKBUF_X2 inst_11361 ( .A(net_9201), .Z(net_11209) );
CLKBUF_X2 inst_13867 ( .A(net_13714), .Z(net_13715) );
AOI22_X2 inst_8158 ( .B1(net_8155), .A1(net_7713), .B2(net_6101), .A2(net_6095), .ZN(net_3994) );
CLKBUF_X2 inst_15080 ( .A(net_14927), .Z(net_14928) );
CLKBUF_X2 inst_12423 ( .A(net_11252), .Z(net_12271) );
NOR2_X2 inst_3461 ( .A1(net_3023), .ZN(net_2756), .A2(net_2498) );
CLKBUF_X2 inst_10974 ( .A(net_9398), .Z(net_10822) );
CLKBUF_X2 inst_9754 ( .A(net_9074), .Z(net_9602) );
MUX2_X2 inst_4969 ( .S(net_2147), .Z(net_1995), .B(net_1994), .A(net_871) );
AOI22_X2 inst_8546 ( .B1(net_6661), .A1(net_6628), .A2(net_6213), .B2(net_6138), .ZN(net_3394) );
CLKBUF_X2 inst_18409 ( .A(net_18256), .Z(net_18257) );
NAND2_X2 inst_4692 ( .ZN(net_2489), .A2(net_2450), .A1(net_2012) );
AOI22_X2 inst_8244 ( .B1(net_8687), .A1(net_8650), .B2(net_6109), .A2(net_3857), .ZN(net_3793) );
NAND2_X2 inst_4883 ( .A2(net_7382), .ZN(net_773), .A1(net_171) );
CLKBUF_X2 inst_10487 ( .A(net_10334), .Z(net_10335) );
AOI22_X2 inst_8580 ( .B1(net_2570), .A2(net_1588), .A1(net_1536), .B2(net_1517), .ZN(net_1514) );
DFFR_X1 inst_7538 ( .Q(net_6478), .D(net_1202), .CK(net_11739), .RN(x6501) );
SDFFR_X2 inst_2178 ( .QN(net_7570), .D(net_3946), .SE(net_3144), .SI(net_2969), .CK(net_10872), .RN(x6501) );
XNOR2_X2 inst_185 ( .A(net_7658), .ZN(net_1646), .B(net_1645) );
CLKBUF_X2 inst_9498 ( .A(net_9345), .Z(net_9346) );
CLKBUF_X2 inst_17474 ( .A(net_17321), .Z(net_17322) );
XNOR2_X2 inst_166 ( .ZN(net_1827), .A(net_1547), .B(net_1540) );
NAND4_X2 inst_3815 ( .ZN(net_3611), .A1(net_3427), .A2(net_3426), .A3(net_3425), .A4(net_3424) );
NAND2_X2 inst_4786 ( .A1(net_2652), .A2(net_2424), .ZN(net_2012) );
CLKBUF_X2 inst_12617 ( .A(net_12464), .Z(net_12465) );
CLKBUF_X2 inst_13822 ( .A(net_13393), .Z(net_13670) );
SDFF_X2 inst_1757 ( .SI(net_7763), .Q(net_7763), .D(net_2711), .SE(net_2560), .CK(net_14248) );
NAND4_X2 inst_3851 ( .ZN(net_1573), .A2(net_1228), .A4(net_1045), .A1(net_744), .A3(net_273) );
INV_X2 inst_6370 ( .ZN(net_1712), .A(net_1711) );
DFF_X1 inst_6772 ( .Q(net_7551), .D(net_4600), .CK(net_12766) );
CLKBUF_X2 inst_12358 ( .A(net_12205), .Z(net_12206) );
CLKBUF_X2 inst_15683 ( .A(net_15530), .Z(net_15531) );
CLKBUF_X2 inst_16143 ( .A(net_15990), .Z(net_15991) );
INV_X2 inst_6359 ( .ZN(net_6056), .A(net_2096) );
CLKBUF_X2 inst_12026 ( .A(net_11873), .Z(net_11874) );
SDFF_X2 inst_1605 ( .Q(net_8114), .D(net_8114), .SI(net_2705), .SE(net_2541), .CK(net_15823) );
CLKBUF_X2 inst_18280 ( .A(net_18127), .Z(net_18128) );
CLKBUF_X2 inst_10206 ( .A(net_10053), .Z(net_10054) );
CLKBUF_X2 inst_11635 ( .A(net_11482), .Z(net_11483) );
CLKBUF_X2 inst_13593 ( .A(net_11020), .Z(net_13441) );
CLKBUF_X2 inst_18518 ( .A(net_18365), .Z(net_18366) );
NAND2_X2 inst_4649 ( .ZN(net_2738), .A2(net_2339), .A1(net_2279) );
CLKBUF_X2 inst_14508 ( .A(net_13014), .Z(net_14356) );
CLKBUF_X2 inst_18462 ( .A(net_18309), .Z(net_18310) );
CLKBUF_X2 inst_12904 ( .A(net_12751), .Z(net_12752) );
CLKBUF_X2 inst_10558 ( .A(net_10405), .Z(net_10406) );
CLKBUF_X2 inst_17975 ( .A(net_15807), .Z(net_17823) );
CLKBUF_X2 inst_12922 ( .A(net_12769), .Z(net_12770) );
CLKBUF_X2 inst_17774 ( .A(net_17621), .Z(net_17622) );
INV_X4 inst_5308 ( .ZN(net_1599), .A(net_1140) );
CLKBUF_X2 inst_15770 ( .A(net_15617), .Z(net_15618) );
CLKBUF_X2 inst_14634 ( .A(net_14481), .Z(net_14482) );
NAND2_X2 inst_4475 ( .ZN(net_4684), .A1(net_4513), .A2(net_4509) );
CLKBUF_X2 inst_17059 ( .A(net_9067), .Z(net_16907) );
AOI22_X2 inst_7757 ( .B1(net_6985), .A1(net_6945), .A2(net_5443), .B2(net_5442), .ZN(net_5378) );
CLKBUF_X2 inst_11077 ( .A(net_10924), .Z(net_10925) );
CLKBUF_X2 inst_16837 ( .A(net_16684), .Z(net_16685) );
CLKBUF_X2 inst_15925 ( .A(net_15772), .Z(net_15773) );
CLKBUF_X2 inst_17514 ( .A(net_17361), .Z(net_17362) );
INV_X4 inst_5201 ( .ZN(net_2863), .A(net_2458) );
CLKBUF_X2 inst_14831 ( .A(net_14678), .Z(net_14679) );
CLKBUF_X2 inst_16121 ( .A(net_15968), .Z(net_15969) );
CLKBUF_X2 inst_16705 ( .A(net_12546), .Z(net_16553) );
SDFFR_X2 inst_2373 ( .SE(net_2260), .Q(net_318), .D(net_318), .CK(net_10460), .RN(x6501), .SI(x3207) );
CLKBUF_X2 inst_11436 ( .A(net_11283), .Z(net_11284) );
CLKBUF_X2 inst_15321 ( .A(net_15168), .Z(net_15169) );
SDFF_X2 inst_1331 ( .Q(net_7946), .D(net_7946), .SE(net_2755), .SI(net_2709), .CK(net_18882) );
CLKBUF_X2 inst_9215 ( .A(net_9062), .Z(net_9063) );
CLKBUF_X2 inst_12322 ( .A(net_12169), .Z(net_12170) );
CLKBUF_X2 inst_15779 ( .A(net_15626), .Z(net_15627) );
DFFR_X1 inst_7404 ( .D(net_5726), .CK(net_13902), .RN(x6501), .Q(x552) );
NOR4_X2 inst_3223 ( .ZN(net_2465), .A4(net_2464), .A2(net_2457), .A3(net_1158), .A1(net_891) );
NOR2_X2 inst_3560 ( .ZN(net_1338), .A1(net_1337), .A2(net_1336) );
SDFFR_X1 inst_2683 ( .SI(net_7546), .SE(net_5043), .CK(net_9692), .RN(x6501), .Q(x3983), .D(x3983) );
CLKBUF_X2 inst_13736 ( .A(net_9519), .Z(net_13584) );
CLKBUF_X2 inst_17442 ( .A(net_17289), .Z(net_17290) );
NAND2_X2 inst_4223 ( .A1(net_6895), .A2(net_5247), .ZN(net_5237) );
CLKBUF_X2 inst_18235 ( .A(net_18082), .Z(net_18083) );
CLKBUF_X2 inst_16910 ( .A(net_16757), .Z(net_16758) );
CLKBUF_X2 inst_14152 ( .A(net_9253), .Z(net_14000) );
CLKBUF_X2 inst_14277 ( .A(net_14124), .Z(net_14125) );
CLKBUF_X2 inst_17182 ( .A(net_17029), .Z(net_17030) );
CLKBUF_X2 inst_13283 ( .A(net_13130), .Z(net_13131) );
HA_X1 inst_6677 ( .S(net_3104), .CO(net_3103), .B(net_2924), .A(x2948) );
CLKBUF_X2 inst_15931 ( .A(net_15778), .Z(net_15779) );
SDFF_X2 inst_1910 ( .D(net_7285), .SI(net_6902), .Q(net_6902), .SE(net_6284), .CK(net_16179) );
CLKBUF_X2 inst_13420 ( .A(net_13267), .Z(net_13268) );
CLKBUF_X2 inst_14461 ( .A(net_9912), .Z(net_14309) );
CLKBUF_X2 inst_16091 ( .A(net_15114), .Z(net_15939) );
CLKBUF_X2 inst_10272 ( .A(net_10119), .Z(net_10120) );
CLKBUF_X2 inst_9265 ( .A(net_9067), .Z(net_9113) );
OAI21_X2 inst_3115 ( .ZN(net_2426), .A(net_2323), .B2(net_2292), .B1(net_2287) );
INV_X4 inst_5814 ( .A(net_7375), .ZN(net_930) );
CLKBUF_X2 inst_15887 ( .A(net_14548), .Z(net_15735) );
NOR4_X2 inst_3219 ( .A1(net_2963), .ZN(net_2779), .A2(net_1841), .A4(net_1115), .A3(net_1041) );
CLKBUF_X2 inst_10867 ( .A(net_9098), .Z(net_10715) );
INV_X4 inst_5673 ( .A(net_7650), .ZN(net_3600) );
CLKBUF_X2 inst_10025 ( .A(net_9347), .Z(net_9873) );
CLKBUF_X2 inst_18659 ( .A(net_18362), .Z(net_18507) );
SDFF_X2 inst_1991 ( .D(net_7266), .SI(net_6843), .Q(net_6843), .SE(net_6282), .CK(net_14310) );
CLKBUF_X2 inst_14872 ( .A(net_9328), .Z(net_14720) );
CLKBUF_X2 inst_13054 ( .A(net_12901), .Z(net_12902) );
OAI21_X2 inst_3066 ( .B2(net_8230), .B1(net_4928), .ZN(net_4724), .A(net_3310) );
AOI22_X2 inst_7861 ( .B2(net_5609), .A2(net_5267), .ZN(net_4580), .B1(net_375), .A1(net_179) );
CLKBUF_X2 inst_14129 ( .A(net_13976), .Z(net_13977) );
CLKBUF_X2 inst_15441 ( .A(net_15288), .Z(net_15289) );
CLKBUF_X2 inst_11630 ( .A(net_11477), .Z(net_11478) );
DFFR_X1 inst_7419 ( .D(net_5532), .CK(net_16620), .RN(x6501), .Q(x653) );
DFF_X1 inst_6771 ( .Q(net_7550), .D(net_4601), .CK(net_12767) );
NAND2_X2 inst_4703 ( .ZN(net_2719), .A2(net_1586), .A1(net_1026) );
INV_X16 inst_6640 ( .ZN(net_3982), .A(net_3327) );
AOI22_X2 inst_8173 ( .B1(net_8862), .A1(net_8307), .B2(net_6252), .A2(net_4345), .ZN(net_3856) );
SDFFR_X1 inst_2672 ( .D(net_6758), .SE(net_4506), .CK(net_11524), .RN(x6501), .SI(x2133), .Q(x2133) );
NOR2_X2 inst_3527 ( .ZN(net_1870), .A2(net_1704), .A1(net_1309) );
CLKBUF_X2 inst_13924 ( .A(net_10202), .Z(net_13772) );
CLKBUF_X2 inst_13637 ( .A(net_13484), .Z(net_13485) );
CLKBUF_X2 inst_9558 ( .A(net_9405), .Z(net_9406) );
INV_X4 inst_6045 ( .A(net_6297), .ZN(net_2640) );
NAND4_X2 inst_3764 ( .ZN(net_4257), .A1(net_3804), .A2(net_3803), .A3(net_3802), .A4(net_3801) );
INV_X2 inst_6408 ( .ZN(net_1068), .A(net_1067) );
AND3_X4 inst_9042 ( .ZN(net_2561), .A3(net_2222), .A1(net_1604), .A2(net_1452) );
AOI221_X2 inst_8764 ( .C2(net_6187), .ZN(net_5464), .B2(net_5463), .A(net_4943), .B1(net_437), .C1(net_200) );
CLKBUF_X2 inst_11912 ( .A(net_11759), .Z(net_11760) );
DFFR_X2 inst_7330 ( .D(net_7643), .QN(net_7640), .CK(net_15643), .RN(x6501) );
CLKBUF_X2 inst_13101 ( .A(net_10095), .Z(net_12949) );
DFFR_X1 inst_7581 ( .Q(net_297), .D(net_274), .CK(net_16322), .RN(x6501) );
SDFFR_X2 inst_2340 ( .SE(net_2757), .D(net_2736), .SI(net_454), .Q(net_454), .CK(net_13854), .RN(x6501) );
CLKBUF_X2 inst_17589 ( .A(net_17436), .Z(net_17437) );
CLKBUF_X2 inst_18324 ( .A(net_15368), .Z(net_18172) );
CLKBUF_X2 inst_15492 ( .A(net_15339), .Z(net_15340) );
CLKBUF_X2 inst_17496 ( .A(net_17343), .Z(net_17344) );
CLKBUF_X2 inst_18027 ( .A(net_17874), .Z(net_17875) );
XOR2_X2 inst_16 ( .Z(net_1426), .B(net_1425), .A(net_707) );
CLKBUF_X2 inst_18562 ( .A(net_18409), .Z(net_18410) );
CLKBUF_X2 inst_15362 ( .A(net_15209), .Z(net_15210) );
CLKBUF_X2 inst_14173 ( .A(net_14020), .Z(net_14021) );
XNOR2_X2 inst_156 ( .ZN(net_1964), .A(net_1963), .B(net_1962) );
OR3_X2 inst_2808 ( .A1(net_6179), .A2(net_6167), .ZN(net_2186), .A3(net_2185) );
CLKBUF_X2 inst_17530 ( .A(net_17377), .Z(net_17378) );
INV_X2 inst_6239 ( .ZN(net_4897), .A(net_4802) );
NOR2_X2 inst_3442 ( .A2(net_3093), .ZN(net_3050), .A1(net_2866) );
SDFFR_X1 inst_2693 ( .SI(net_7555), .SE(net_5043), .CK(net_12735), .RN(x6501), .Q(x3847), .D(x3847) );
CLKBUF_X2 inst_14920 ( .A(net_14767), .Z(net_14768) );
CLKBUF_X2 inst_17228 ( .A(net_14724), .Z(net_17076) );
CLKBUF_X2 inst_10307 ( .A(net_10154), .Z(net_10155) );
CLKBUF_X2 inst_18133 ( .A(net_9996), .Z(net_17981) );
INV_X4 inst_5380 ( .A(net_2093), .ZN(net_1350) );
CLKBUF_X2 inst_14838 ( .A(net_14685), .Z(net_14686) );
CLKBUF_X2 inst_10936 ( .A(net_10783), .Z(net_10784) );
INV_X2 inst_6473 ( .A(net_6794), .ZN(net_844) );
SDFF_X2 inst_1549 ( .Q(net_7978), .D(net_7978), .SI(net_2705), .SE(net_2542), .CK(net_15832) );
OAI21_X2 inst_3020 ( .B2(net_5044), .ZN(net_5040), .A(net_4885), .B1(net_1938) );
INV_X2 inst_6186 ( .ZN(net_5828), .A(net_5779) );
CLKBUF_X2 inst_9239 ( .A(net_9086), .Z(net_9087) );
CLKBUF_X2 inst_12894 ( .A(net_12741), .Z(net_12742) );
CLKBUF_X2 inst_10576 ( .A(net_10423), .Z(net_10424) );
CLKBUF_X2 inst_13477 ( .A(net_13324), .Z(net_13325) );
SDFF_X2 inst_821 ( .SI(net_8513), .Q(net_8513), .D(net_3951), .SE(net_3884), .CK(net_13392) );
OR2_X2 inst_2881 ( .ZN(net_2517), .A2(net_2414), .A1(net_258) );
AND2_X4 inst_9113 ( .A1(net_7217), .ZN(net_6173), .A2(net_1733) );
AOI21_X2 inst_8879 ( .B2(net_5871), .ZN(net_5866), .A(net_5865), .B1(x240) );
CLKBUF_X2 inst_16225 ( .A(net_13585), .Z(net_16073) );
SDFF_X2 inst_980 ( .SI(net_7316), .Q(net_6723), .D(net_6723), .SE(net_3124), .CK(net_9881) );
CLKBUF_X2 inst_15750 ( .A(net_15597), .Z(net_15598) );
CLKBUF_X2 inst_16021 ( .A(net_15868), .Z(net_15869) );
AOI22_X2 inst_8486 ( .B1(net_6677), .A1(net_6644), .A2(net_6213), .B2(net_6138), .ZN(net_3454) );
CLKBUF_X2 inst_16714 ( .A(net_12751), .Z(net_16562) );
SDFF_X2 inst_1785 ( .D(net_7297), .SI(net_6994), .Q(net_6994), .SE(net_6283), .CK(net_18189) );
CLKBUF_X2 inst_10104 ( .A(net_9951), .Z(net_9952) );
CLKBUF_X2 inst_12939 ( .A(net_12786), .Z(net_12787) );
NAND2_X2 inst_4213 ( .A1(net_6890), .ZN(net_5248), .A2(net_5247) );
CLKBUF_X2 inst_9341 ( .A(net_9099), .Z(net_9189) );
CLKBUF_X2 inst_15180 ( .A(net_10987), .Z(net_15028) );
CLKBUF_X2 inst_9575 ( .A(net_9422), .Z(net_9423) );
SDFFR_X2 inst_2286 ( .SE(net_2801), .D(net_1330), .SI(net_204), .Q(net_204), .CK(net_14960), .RN(x6501) );
INV_X4 inst_6022 ( .A(net_7652), .ZN(net_1568) );
CLKBUF_X2 inst_10694 ( .A(net_10541), .Z(net_10542) );
CLKBUF_X2 inst_12118 ( .A(net_11965), .Z(net_11966) );
CLKBUF_X2 inst_19158 ( .A(net_19005), .Z(net_19006) );
DFFR_X2 inst_7142 ( .QN(net_9056), .D(net_2966), .CK(net_11160), .RN(x6501) );
DFFR_X1 inst_7512 ( .D(net_1434), .Q(net_280), .CK(net_16611), .RN(x6501) );
SDFFR_X2 inst_2137 ( .SI(net_7177), .Q(net_7177), .D(net_6428), .SE(net_4362), .CK(net_13726), .RN(x6501) );
CLKBUF_X2 inst_9406 ( .A(net_9253), .Z(net_9254) );
DFFR_X2 inst_7107 ( .QN(net_6333), .D(net_3188), .CK(net_18961), .RN(x6501) );
SDFF_X2 inst_1613 ( .Q(net_8120), .D(net_8120), .SI(net_2702), .SE(net_2541), .CK(net_18038) );
INV_X16 inst_6624 ( .ZN(net_4190), .A(net_3571) );
CLKBUF_X2 inst_16503 ( .A(net_16350), .Z(net_16351) );
INV_X4 inst_5659 ( .A(net_7395), .ZN(net_939) );
CLKBUF_X2 inst_15508 ( .A(net_15323), .Z(net_15356) );
INV_X4 inst_5965 ( .A(net_6402), .ZN(net_2810) );
CLKBUF_X2 inst_15098 ( .A(net_14945), .Z(net_14946) );
CLKBUF_X2 inst_17002 ( .A(net_16849), .Z(net_16850) );
SDFF_X2 inst_1141 ( .SI(net_7311), .Q(net_6586), .D(net_6586), .SE(net_3069), .CK(net_9906) );
CLKBUF_X2 inst_15982 ( .A(net_15708), .Z(net_15830) );
SDFFR_X2 inst_2488 ( .D(net_7366), .SE(net_2548), .SI(net_2546), .QN(net_259), .CK(net_13543), .RN(x6501) );
NOR2_X2 inst_3589 ( .A1(net_7518), .ZN(net_1336), .A2(net_538) );
CLKBUF_X2 inst_18379 ( .A(net_18226), .Z(net_18227) );
SDFF_X2 inst_932 ( .SI(net_7340), .Q(net_6681), .D(net_6681), .SE(net_3126), .CK(net_9509) );
XNOR2_X2 inst_180 ( .B(net_4697), .ZN(net_1676), .A(net_1321) );
CLKBUF_X2 inst_12891 ( .A(net_12738), .Z(net_12739) );
CLKBUF_X2 inst_13472 ( .A(net_9842), .Z(net_13320) );
AND2_X4 inst_9057 ( .ZN(net_3329), .A1(net_3328), .A2(net_3325) );
CLKBUF_X2 inst_18762 ( .A(net_18609), .Z(net_18610) );
CLKBUF_X2 inst_16584 ( .A(net_10586), .Z(net_16432) );
AOI22_X2 inst_8003 ( .B1(net_8079), .A1(net_7739), .B2(net_6108), .A2(net_6096), .ZN(net_4131) );
CLKBUF_X2 inst_15474 ( .A(net_15321), .Z(net_15322) );
AOI22_X2 inst_8475 ( .B1(net_6608), .A1(net_6575), .A2(net_6257), .B2(net_6110), .ZN(net_3465) );
CLKBUF_X2 inst_11995 ( .A(net_11842), .Z(net_11843) );
INV_X2 inst_6455 ( .A(net_8967), .ZN(net_587) );
CLKBUF_X2 inst_12635 ( .A(net_12482), .Z(net_12483) );
CLKBUF_X2 inst_12654 ( .A(net_12501), .Z(net_12502) );
CLKBUF_X2 inst_17870 ( .A(net_17717), .Z(net_17718) );
CLKBUF_X2 inst_10318 ( .A(net_9570), .Z(net_10166) );
CLKBUF_X2 inst_13527 ( .A(net_13374), .Z(net_13375) );
CLKBUF_X2 inst_15214 ( .A(net_13234), .Z(net_15062) );
NOR3_X2 inst_3287 ( .ZN(net_6264), .A3(net_6251), .A1(net_6179), .A2(net_3161) );
XNOR2_X2 inst_211 ( .ZN(net_1463), .A(net_1462), .B(net_823) );
INV_X4 inst_5892 ( .A(net_8290), .ZN(net_1243) );
CLKBUF_X2 inst_11628 ( .A(net_9985), .Z(net_11476) );
NAND2_X2 inst_4659 ( .ZN(net_2266), .A1(net_2262), .A2(net_2078) );
OAI21_X2 inst_3120 ( .ZN(net_2294), .A(net_2293), .B2(net_2292), .B1(net_2224) );
INV_X4 inst_5735 ( .A(net_7523), .ZN(net_625) );
INV_X4 inst_5917 ( .A(net_7577), .ZN(net_529) );
CLKBUF_X2 inst_18579 ( .A(net_18426), .Z(net_18427) );
CLKBUF_X2 inst_18934 ( .A(net_18781), .Z(net_18782) );
CLKBUF_X2 inst_11565 ( .A(net_11412), .Z(net_11413) );
CLKBUF_X2 inst_15243 ( .A(net_15090), .Z(net_15091) );
CLKBUF_X2 inst_17004 ( .A(net_16851), .Z(net_16852) );
DFFS_X1 inst_6945 ( .D(net_6145), .CK(net_13633), .SN(x6501), .Q(x771) );
CLKBUF_X2 inst_12806 ( .A(net_12653), .Z(net_12654) );
SDFFR_X1 inst_2736 ( .SI(net_9049), .Q(net_9049), .SE(net_3208), .D(net_3127), .CK(net_10650), .RN(x6501) );
DFFR_X2 inst_7178 ( .QN(net_8904), .D(net_2516), .CK(net_16297), .RN(x6501) );
CLKBUF_X2 inst_18138 ( .A(net_17985), .Z(net_17986) );
NAND2_X2 inst_4489 ( .A1(net_7198), .A2(net_5655), .ZN(net_4483) );
CLKBUF_X2 inst_17015 ( .A(net_16862), .Z(net_16863) );
INV_X4 inst_5523 ( .A(net_956), .ZN(net_668) );
CLKBUF_X2 inst_10637 ( .A(net_10484), .Z(net_10485) );
SDFF_X2 inst_1403 ( .Q(net_8183), .D(net_8183), .SI(net_2655), .SE(net_2561), .CK(net_15460) );
DFFR_X2 inst_7155 ( .QN(net_5949), .D(net_2853), .CK(net_11152), .RN(x6501) );
CLKBUF_X2 inst_14811 ( .A(net_12475), .Z(net_14659) );
CLKBUF_X2 inst_15100 ( .A(net_14947), .Z(net_14948) );
CLKBUF_X2 inst_14684 ( .A(net_14531), .Z(net_14532) );
CLKBUF_X2 inst_18745 ( .A(net_18592), .Z(net_18593) );
XOR2_X2 inst_42 ( .Z(net_1045), .A(net_654), .B(net_190) );
CLKBUF_X2 inst_10521 ( .A(net_9298), .Z(net_10369) );
CLKBUF_X2 inst_13535 ( .A(net_9353), .Z(net_13383) );
CLKBUF_X2 inst_15880 ( .A(net_15727), .Z(net_15728) );
CLKBUF_X2 inst_16009 ( .A(net_13334), .Z(net_15857) );
CLKBUF_X2 inst_17732 ( .A(net_17579), .Z(net_17580) );
NAND2_X2 inst_4084 ( .A1(net_7623), .A2(net_5751), .ZN(net_5750) );
CLKBUF_X2 inst_16154 ( .A(net_16001), .Z(net_16002) );
SDFF_X2 inst_1479 ( .SI(net_7292), .Q(net_7069), .D(net_7069), .SE(net_6280), .CK(net_14919) );
CLKBUF_X2 inst_18346 ( .A(net_18193), .Z(net_18194) );
SDFF_X2 inst_437 ( .Q(net_8765), .D(net_8765), .SE(net_3982), .SI(net_3955), .CK(net_13282) );
CLKBUF_X2 inst_11606 ( .A(net_11453), .Z(net_11454) );
CLKBUF_X2 inst_16664 ( .A(net_15296), .Z(net_16512) );
CLKBUF_X2 inst_13307 ( .A(net_13154), .Z(net_13155) );
AOI22_X2 inst_8316 ( .B1(net_8558), .A1(net_8447), .A2(net_6263), .B2(net_6262), .ZN(net_3729) );
CLKBUF_X2 inst_14489 ( .A(net_14336), .Z(net_14337) );
CLKBUF_X2 inst_14391 ( .A(net_14238), .Z(net_14239) );
CLKBUF_X2 inst_16034 ( .A(net_9794), .Z(net_15882) );
CLKBUF_X2 inst_17513 ( .A(net_17360), .Z(net_17361) );
CLKBUF_X2 inst_12782 ( .A(net_9332), .Z(net_12630) );
CLKBUF_X2 inst_9425 ( .A(net_9272), .Z(net_9273) );
CLKBUF_X2 inst_10451 ( .A(net_9635), .Z(net_10299) );
SDFF_X2 inst_1706 ( .Q(net_7891), .D(net_7891), .SI(net_2719), .SE(net_2543), .CK(net_15963) );
DFF_X1 inst_6733 ( .Q(net_6778), .D(net_5636), .CK(net_9207) );
DFF_X1 inst_6778 ( .Q(net_7529), .D(net_4594), .CK(net_9541) );
CLKBUF_X2 inst_17638 ( .A(net_12124), .Z(net_17486) );
SDFFR_X2 inst_2220 ( .Q(net_7456), .D(net_7456), .SE(net_2863), .CK(net_10631), .SI(x13534), .RN(x6501) );
CLKBUF_X2 inst_18769 ( .A(net_18616), .Z(net_18617) );
CLKBUF_X2 inst_17075 ( .A(net_16922), .Z(net_16923) );
CLKBUF_X2 inst_9958 ( .A(net_9805), .Z(net_9806) );
SDFFR_X2 inst_2247 ( .SE(net_5582), .D(net_2637), .CK(net_14203), .RN(x6501), .SI(x132), .Q(x132) );
CLKBUF_X2 inst_13517 ( .A(net_13364), .Z(net_13365) );
CLKBUF_X2 inst_9706 ( .A(net_9553), .Z(net_9554) );
CLKBUF_X2 inst_11852 ( .A(net_11699), .Z(net_11700) );
CLKBUF_X2 inst_17302 ( .A(net_17149), .Z(net_17150) );
INV_X4 inst_5786 ( .A(net_6361), .ZN(net_690) );
NOR2_X2 inst_3418 ( .ZN(net_3249), .A1(net_3177), .A2(net_3176) );
CLKBUF_X2 inst_17784 ( .A(net_17631), .Z(net_17632) );
NOR2_X4 inst_3334 ( .ZN(net_2321), .A1(net_2170), .A2(net_777) );
SDFF_X2 inst_407 ( .SI(net_8321), .Q(net_8321), .SE(net_3978), .D(net_3955), .CK(net_11023) );
NOR2_X2 inst_3558 ( .ZN(net_3038), .A2(net_1345), .A1(net_561) );
SDFF_X2 inst_1208 ( .Q(net_7973), .D(net_7973), .SE(net_2755), .SI(net_2716), .CK(net_17109) );
INV_X4 inst_5843 ( .A(net_7174), .ZN(net_2957) );
SDFF_X2 inst_652 ( .Q(net_8424), .D(net_8424), .SI(net_3944), .SE(net_3934), .CK(net_10835) );
CLKBUF_X2 inst_15643 ( .A(net_15490), .Z(net_15491) );
CLKBUF_X2 inst_9935 ( .A(net_9552), .Z(net_9783) );
SDFF_X2 inst_677 ( .Q(net_8696), .D(net_8696), .SI(net_3952), .SE(net_3935), .CK(net_12880) );
XNOR2_X2 inst_130 ( .ZN(net_2824), .A(net_2550), .B(net_807) );
CLKBUF_X2 inst_12155 ( .A(net_10029), .Z(net_12003) );
SDFF_X2 inst_1566 ( .Q(net_8040), .D(net_8040), .SI(net_2704), .SE(net_2545), .CK(net_16996) );
CLKBUF_X2 inst_12468 ( .A(net_12315), .Z(net_12316) );
CLKBUF_X2 inst_10829 ( .A(net_9901), .Z(net_10677) );
CLKBUF_X2 inst_14892 ( .A(net_14739), .Z(net_14740) );
CLKBUF_X2 inst_10489 ( .A(net_10336), .Z(net_10337) );
CLKBUF_X2 inst_18247 ( .A(net_18094), .Z(net_18095) );
SDFF_X2 inst_1054 ( .SI(net_7325), .Q(net_6666), .D(net_6666), .SE(net_3126), .CK(net_11329) );
CLKBUF_X2 inst_18650 ( .A(net_18497), .Z(net_18498) );
CLKBUF_X2 inst_11420 ( .A(net_11267), .Z(net_11268) );
SDFF_X2 inst_972 ( .SI(net_7335), .Q(net_6742), .D(net_6742), .SE(net_3124), .CK(net_9769) );
CLKBUF_X2 inst_15227 ( .A(net_15074), .Z(net_15075) );
CLKBUF_X2 inst_13992 ( .A(net_13839), .Z(net_13840) );
SDFF_X2 inst_1843 ( .D(net_7284), .SI(net_7021), .Q(net_7021), .SE(net_6277), .CK(net_16193) );
CLKBUF_X2 inst_16897 ( .A(net_16744), .Z(net_16745) );
CLKBUF_X2 inst_16639 ( .A(net_16486), .Z(net_16487) );
CLKBUF_X2 inst_11113 ( .A(net_10668), .Z(net_10961) );
CLKBUF_X2 inst_18853 ( .A(net_11114), .Z(net_18701) );
CLKBUF_X2 inst_10224 ( .A(net_10071), .Z(net_10072) );
CLKBUF_X2 inst_11951 ( .A(net_11798), .Z(net_11799) );
CLKBUF_X2 inst_11480 ( .A(net_11327), .Z(net_11328) );
CLKBUF_X2 inst_14679 ( .A(net_14526), .Z(net_14527) );
CLKBUF_X2 inst_15392 ( .A(net_15239), .Z(net_15240) );
CLKBUF_X2 inst_12717 ( .A(net_12564), .Z(net_12565) );
XNOR2_X2 inst_204 ( .ZN(net_1539), .B(net_1201), .A(net_1194) );
SDFF_X2 inst_1550 ( .Q(net_8006), .D(net_8006), .SI(net_2704), .SE(net_2542), .CK(net_17004) );
SDFF_X2 inst_910 ( .SI(net_8729), .Q(net_8729), .SE(net_6195), .D(net_3954), .CK(net_10885) );
CLKBUF_X2 inst_14816 ( .A(net_10302), .Z(net_14664) );
CLKBUF_X2 inst_10134 ( .A(net_9556), .Z(net_9982) );
AOI221_X2 inst_8772 ( .B2(net_8239), .ZN(net_5269), .B1(net_5268), .C2(net_5267), .A(net_4917), .C1(net_176) );
CLKBUF_X2 inst_13080 ( .A(net_12927), .Z(net_12928) );
CLKBUF_X2 inst_16207 ( .A(net_16054), .Z(net_16055) );
CLKBUF_X2 inst_12494 ( .A(net_12341), .Z(net_12342) );
DFFR_X1 inst_7562 ( .Q(net_6415), .D(net_6412), .CK(net_9663), .RN(x6501) );
CLKBUF_X2 inst_12344 ( .A(net_12191), .Z(net_12192) );
CLKBUF_X2 inst_11515 ( .A(net_11362), .Z(net_11363) );
SDFF_X2 inst_937 ( .SI(net_7315), .Q(net_6656), .D(net_6656), .SE(net_3126), .CK(net_9955) );
DFFR_X1 inst_7401 ( .D(net_5742), .CK(net_14051), .RN(x6501), .Q(x258) );
CLKBUF_X2 inst_15315 ( .A(net_15162), .Z(net_15163) );
SDFF_X2 inst_355 ( .Q(net_8743), .D(net_8743), .SE(net_3982), .SI(net_3980), .CK(net_10748) );
CLKBUF_X2 inst_9259 ( .A(net_9106), .Z(net_9107) );
INV_X2 inst_6584 ( .A(net_7167), .ZN(net_478) );
NOR2_X2 inst_3498 ( .ZN(net_1937), .A1(net_1936), .A2(net_1935) );
DFF_X1 inst_6753 ( .Q(net_6763), .D(net_5613), .CK(net_10488) );
CLKBUF_X2 inst_16139 ( .A(net_14528), .Z(net_15987) );
NAND4_X2 inst_3693 ( .ZN(net_4444), .A4(net_4344), .A1(net_3807), .A2(net_3806), .A3(net_3805) );
DFF_X1 inst_6806 ( .Q(net_8223), .D(net_4422), .CK(net_16556) );
CLKBUF_X2 inst_11309 ( .A(net_11156), .Z(net_11157) );
CLKBUF_X2 inst_14619 ( .A(net_14466), .Z(net_14467) );
CLKBUF_X2 inst_15655 ( .A(net_15502), .Z(net_15503) );
CLKBUF_X2 inst_18614 ( .A(net_17627), .Z(net_18462) );
NAND4_X2 inst_3769 ( .ZN(net_4252), .A1(net_3772), .A2(net_3771), .A3(net_3770), .A4(net_3769) );
NAND2_X4 inst_4053 ( .A2(net_8902), .ZN(net_6123), .A1(net_1724) );
CLKBUF_X2 inst_16466 ( .A(net_16313), .Z(net_16314) );
SDFF_X2 inst_1747 ( .Q(net_8212), .D(net_8212), .SI(net_2656), .SE(net_2561), .CK(net_16706) );
INV_X4 inst_5109 ( .ZN(net_4947), .A(net_4880) );
AND2_X4 inst_9066 ( .ZN(net_6137), .A2(net_3248), .A1(net_3247) );
CLKBUF_X2 inst_10477 ( .A(net_10324), .Z(net_10325) );
CLKBUF_X2 inst_11834 ( .A(net_9136), .Z(net_11682) );
CLKBUF_X2 inst_11978 ( .A(net_11825), .Z(net_11826) );
CLKBUF_X2 inst_13026 ( .A(net_12873), .Z(net_12874) );
CLKBUF_X2 inst_13352 ( .A(net_13199), .Z(net_13200) );
NAND3_X2 inst_3917 ( .ZN(net_5621), .A1(net_5550), .A3(net_5484), .A2(net_5323) );
CLKBUF_X2 inst_9419 ( .A(net_9266), .Z(net_9267) );
CLKBUF_X2 inst_13243 ( .A(net_9610), .Z(net_13091) );
SDFFR_X2 inst_2574 ( .QN(net_6379), .SE(net_2147), .D(net_2041), .SI(net_1947), .CK(net_18126), .RN(x6501) );
SDFFR_X2 inst_2229 ( .Q(net_7471), .D(net_7471), .SE(net_2863), .CK(net_12174), .SI(x13423), .RN(x6501) );
CLKBUF_X2 inst_11456 ( .A(net_11303), .Z(net_11304) );
CLKBUF_X2 inst_16613 ( .A(net_16460), .Z(net_16461) );
CLKBUF_X2 inst_16966 ( .A(net_16813), .Z(net_16814) );
INV_X2 inst_6252 ( .ZN(net_4852), .A(net_4738) );
CLKBUF_X2 inst_14587 ( .A(net_14434), .Z(net_14435) );
SDFF_X2 inst_1245 ( .SI(net_7687), .Q(net_7687), .D(net_2719), .SE(net_2714), .CK(net_18821) );
CLKBUF_X2 inst_19131 ( .A(net_16230), .Z(net_18979) );
CLKBUF_X2 inst_12560 ( .A(net_9192), .Z(net_12408) );
CLKBUF_X2 inst_16941 ( .A(net_16788), .Z(net_16789) );
NAND4_X2 inst_3788 ( .ZN(net_4233), .A1(net_3653), .A2(net_3652), .A3(net_3651), .A4(net_3650) );
INV_X4 inst_5409 ( .A(net_1480), .ZN(net_1138) );
NAND4_X2 inst_3663 ( .A4(net_6016), .A1(net_6015), .ZN(net_4602), .A2(net_4114), .A3(net_4113) );
CLKBUF_X2 inst_11977 ( .A(net_11824), .Z(net_11825) );
CLKBUF_X2 inst_15526 ( .A(net_15373), .Z(net_15374) );
OAI21_X2 inst_3008 ( .B2(net_5755), .ZN(net_5741), .A(net_5740), .B1(net_631) );
INV_X4 inst_5515 ( .ZN(net_882), .A(net_771) );
INV_X4 inst_5900 ( .A(net_9013), .ZN(net_894) );
AOI22_X2 inst_8234 ( .B1(net_8575), .A1(net_8464), .A2(net_6263), .B2(net_6262), .ZN(net_3803) );
CLKBUF_X2 inst_10640 ( .A(net_10487), .Z(net_10488) );
NAND2_X2 inst_4071 ( .A2(net_6788), .ZN(net_5776), .A1(net_5775) );
AOI221_X4 inst_8738 ( .B1(net_8712), .C1(net_8490), .B2(net_4350), .C2(net_4349), .ZN(net_4328), .A(net_4232) );
CLKBUF_X2 inst_13614 ( .A(net_13461), .Z(net_13462) );
CLKBUF_X2 inst_11363 ( .A(net_11210), .Z(net_11211) );
AOI22_X2 inst_8249 ( .B1(net_8799), .A1(net_8540), .ZN(net_6224), .A2(net_3861), .B2(net_3860) );
SDFFR_X2 inst_2469 ( .D(net_6318), .SE(net_2678), .SI(net_440), .Q(net_440), .CK(net_17445), .RN(x6501) );
AOI22_X2 inst_7868 ( .B2(net_5609), .A2(net_5267), .ZN(net_4573), .B1(net_359), .A1(net_163) );
CLKBUF_X2 inst_9287 ( .A(net_9134), .Z(net_9135) );
CLKBUF_X2 inst_13230 ( .A(net_10747), .Z(net_13078) );
NAND2_X2 inst_4736 ( .ZN(net_2710), .A1(net_1650), .A2(net_1586) );
CLKBUF_X2 inst_16509 ( .A(net_16356), .Z(net_16357) );
AOI22_X2 inst_8437 ( .B1(net_6732), .A1(net_6699), .B2(net_6202), .A2(net_3520), .ZN(net_3504) );
CLKBUF_X2 inst_14442 ( .A(net_11065), .Z(net_14290) );
CLKBUF_X2 inst_14761 ( .A(net_14608), .Z(net_14609) );
INV_X2 inst_6259 ( .ZN(net_4639), .A(net_4547) );
CLKBUF_X2 inst_17417 ( .A(net_16622), .Z(net_17265) );
CLKBUF_X2 inst_10330 ( .A(net_9938), .Z(net_10178) );
NAND4_X2 inst_3715 ( .ZN(net_4422), .A4(net_4329), .A1(net_3666), .A2(net_3665), .A3(net_3664) );
DFFR_X2 inst_6983 ( .QN(net_5959), .D(net_5897), .CK(net_11495), .RN(x6501) );
CLKBUF_X2 inst_10929 ( .A(net_10776), .Z(net_10777) );
CLKBUF_X2 inst_16733 ( .A(net_16580), .Z(net_16581) );
OAI21_X2 inst_3042 ( .B2(net_8245), .B1(net_4928), .ZN(net_4808), .A(net_3385) );
CLKBUF_X2 inst_17328 ( .A(net_14322), .Z(net_17176) );
SDFF_X2 inst_981 ( .SI(net_7317), .Q(net_6724), .D(net_6724), .SE(net_3124), .CK(net_9879) );
AOI22_X4 inst_7735 ( .B1(net_8188), .A1(net_7678), .B2(net_6099), .A2(net_4399), .ZN(net_3999) );
CLKBUF_X2 inst_11940 ( .A(net_11787), .Z(net_11788) );
AOI221_X2 inst_8815 ( .C2(net_5535), .B2(net_5260), .A(net_4898), .ZN(net_4712), .B1(net_3051), .C1(net_458) );
CLKBUF_X2 inst_17746 ( .A(net_15479), .Z(net_17594) );
INV_X2 inst_6189 ( .ZN(net_5787), .A(net_5753) );
CLKBUF_X2 inst_12260 ( .A(net_10057), .Z(net_12108) );
CLKBUF_X2 inst_12064 ( .A(net_10065), .Z(net_11912) );
CLKBUF_X2 inst_15056 ( .A(net_13849), .Z(net_14904) );
SDFFS_X2 inst_2094 ( .SI(net_7261), .Q(net_6382), .D(net_6382), .SE(net_2147), .CK(net_15015), .SN(x6501) );
NOR2_X2 inst_3417 ( .ZN(net_3373), .A1(net_3180), .A2(net_3179) );
INV_X2 inst_6279 ( .ZN(net_4230), .A(net_4213) );
DFF_X1 inst_6794 ( .QN(net_8241), .D(net_4439), .CK(net_17600) );
CLKBUF_X2 inst_13347 ( .A(net_13121), .Z(net_13195) );
INV_X4 inst_5406 ( .ZN(net_1673), .A(net_876) );
CLKBUF_X2 inst_14337 ( .A(net_14184), .Z(net_14185) );
INV_X2 inst_6292 ( .ZN(net_4206), .A(net_3915) );
CLKBUF_X2 inst_14947 ( .A(net_12622), .Z(net_14795) );
CLKBUF_X2 inst_13959 ( .A(net_13806), .Z(net_13807) );
INV_X4 inst_5324 ( .ZN(net_5691), .A(net_1366) );
NOR2_X2 inst_3491 ( .A1(net_2652), .ZN(net_2308), .A2(net_2161) );
SDFFR_X2 inst_2393 ( .SE(net_2260), .Q(net_360), .D(net_360), .CK(net_10406), .RN(x6501), .SI(x1935) );
XOR2_X1 inst_71 ( .Z(net_3541), .A(net_3267), .B(x2856) );
CLKBUF_X2 inst_14787 ( .A(net_14634), .Z(net_14635) );
NAND2_X2 inst_4079 ( .A2(net_6784), .A1(net_5835), .ZN(net_5767) );
CLKBUF_X2 inst_10114 ( .A(net_9961), .Z(net_9962) );
NOR4_X2 inst_3231 ( .ZN(net_2083), .A3(net_1795), .A2(net_1793), .A4(net_1791), .A1(net_1789) );
AND2_X4 inst_9084 ( .ZN(net_2776), .A2(net_2775), .A1(net_1564) );
CLKBUF_X2 inst_16902 ( .A(net_16749), .Z(net_16750) );
CLKBUF_X2 inst_12884 ( .A(net_12731), .Z(net_12732) );
CLKBUF_X2 inst_14407 ( .A(net_14254), .Z(net_14255) );
CLKBUF_X2 inst_16833 ( .A(net_16680), .Z(net_16681) );
XNOR2_X2 inst_336 ( .B(net_7375), .A(net_6357), .ZN(net_786) );
CLKBUF_X2 inst_12129 ( .A(net_11976), .Z(net_11977) );
CLKBUF_X2 inst_16923 ( .A(net_16770), .Z(net_16771) );
INV_X2 inst_6479 ( .ZN(net_900), .A(net_209) );
SDFF_X2 inst_1939 ( .SI(net_8073), .Q(net_8073), .D(net_2660), .SE(net_2508), .CK(net_16975) );
INV_X4 inst_5157 ( .A(net_3152), .ZN(net_3151) );
CLKBUF_X2 inst_18872 ( .A(net_18142), .Z(net_18720) );
OAI33_X1 inst_2902 ( .B1(net_4924), .ZN(net_4822), .A2(net_4821), .B3(net_4685), .A3(net_4474), .B2(net_2255), .A1(net_2098) );
CLKBUF_X2 inst_14503 ( .A(net_14350), .Z(net_14351) );
AOI22_X2 inst_7844 ( .A1(net_7180), .A2(net_5655), .B2(net_5520), .ZN(net_4664), .B1(net_287) );
CLKBUF_X2 inst_17424 ( .A(net_12310), .Z(net_17272) );
AOI221_X4 inst_8726 ( .B1(net_8729), .C1(net_8507), .B2(net_4350), .C2(net_4349), .ZN(net_4339), .A(net_4250) );
INV_X4 inst_5174 ( .ZN(net_3087), .A(net_2961) );
AOI22_X2 inst_8508 ( .B1(net_6522), .A1(net_6489), .A2(net_6137), .B2(net_6104), .ZN(net_3432) );
CLKBUF_X2 inst_9553 ( .A(net_9400), .Z(net_9401) );
CLKBUF_X2 inst_13450 ( .A(net_10538), .Z(net_13298) );
CLKBUF_X2 inst_11736 ( .A(net_11459), .Z(net_11584) );
AOI22_X2 inst_8263 ( .B1(net_8727), .A1(net_8505), .B2(net_4350), .A2(net_4349), .ZN(net_3775) );
INV_X4 inst_5870 ( .A(net_7250), .ZN(net_1944) );
CLKBUF_X2 inst_17218 ( .A(net_14032), .Z(net_17066) );
INV_X4 inst_5998 ( .A(net_6347), .ZN(net_2739) );
CLKBUF_X2 inst_18432 ( .A(net_18279), .Z(net_18280) );
CLKBUF_X2 inst_17352 ( .A(net_17199), .Z(net_17200) );
CLKBUF_X2 inst_18593 ( .A(net_15736), .Z(net_18441) );
NAND4_X2 inst_3752 ( .ZN(net_4278), .A1(net_4002), .A2(net_4001), .A3(net_4000), .A4(net_3999) );
XNOR2_X2 inst_284 ( .A(net_1780), .ZN(net_1013), .B(net_202) );
CLKBUF_X2 inst_13809 ( .A(net_13656), .Z(net_13657) );
CLKBUF_X2 inst_16756 ( .A(net_16603), .Z(net_16604) );
SDFFR_X2 inst_2579 ( .D(net_7387), .QN(net_7247), .SI(net_1957), .SE(net_1379), .CK(net_18116), .RN(x6501) );
SDFF_X2 inst_1713 ( .Q(net_7980), .D(net_7980), .SI(net_2709), .SE(net_2542), .CK(net_15746) );
CLKBUF_X2 inst_12668 ( .A(net_9638), .Z(net_12516) );
INV_X4 inst_5650 ( .A(net_7230), .ZN(net_1810) );
DFFR_X2 inst_6970 ( .QN(net_6285), .D(net_5928), .CK(net_13884), .RN(x6501) );
NAND2_X2 inst_4527 ( .A2(net_3566), .ZN(net_3559), .A1(net_3555) );
CLKBUF_X2 inst_9532 ( .A(net_9379), .Z(net_9380) );
OAI21_X2 inst_3137 ( .B2(net_2063), .ZN(net_2062), .A(net_2056), .B1(net_734) );
CLKBUF_X2 inst_16632 ( .A(net_9415), .Z(net_16480) );
CLKBUF_X2 inst_11668 ( .A(net_11515), .Z(net_11516) );
CLKBUF_X2 inst_18337 ( .A(net_18184), .Z(net_18185) );
INV_X4 inst_5437 ( .ZN(net_1962), .A(net_1175) );
DFFR_X1 inst_7544 ( .D(net_1052), .Q(net_295), .CK(net_11635), .RN(x6501) );
NAND2_X2 inst_4496 ( .ZN(net_4476), .A2(net_4388), .A1(net_2620) );
DFFR_X2 inst_7357 ( .Q(net_7335), .CK(net_9437), .D(x12962), .RN(x6501) );
INV_X2 inst_6344 ( .ZN(net_2446), .A(net_2445) );
SDFF_X2 inst_951 ( .SI(net_7336), .Q(net_6710), .D(net_6710), .SE(net_3125), .CK(net_9507) );
CLKBUF_X2 inst_12565 ( .A(net_12412), .Z(net_12413) );
CLKBUF_X1 inst_7727 ( .A(x192486), .Z(x999) );
CLKBUF_X2 inst_9836 ( .A(net_9547), .Z(net_9684) );
INV_X4 inst_5831 ( .A(net_8260), .ZN(net_2997) );
CLKBUF_X2 inst_15414 ( .A(net_13593), .Z(net_15262) );
CLKBUF_X2 inst_10268 ( .A(net_9147), .Z(net_10116) );
CLKBUF_X2 inst_11253 ( .A(net_10285), .Z(net_11101) );
AOI21_X2 inst_8938 ( .B2(net_5784), .ZN(net_5663), .A(net_5659), .B1(x394) );
OAI211_X2 inst_3188 ( .C2(net_6444), .C1(net_4950), .ZN(net_4823), .A(net_4652), .B(net_4498) );
DFFR_X2 inst_7358 ( .Q(net_7326), .CK(net_11762), .D(x13038), .RN(x6501) );
DFFR_X2 inst_7351 ( .Q(net_7315), .CK(net_11378), .D(x13145), .RN(x6501) );
DFFR_X1 inst_7435 ( .QN(net_8915), .D(net_4851), .CK(net_16692), .RN(x6501) );
CLKBUF_X2 inst_11545 ( .A(net_11295), .Z(net_11393) );
OAI21_X2 inst_3129 ( .A(net_5951), .B2(net_2849), .ZN(net_2209), .B1(net_1732) );
NAND2_X2 inst_4674 ( .ZN(net_2378), .A1(net_2115), .A2(net_2113) );
CLKBUF_X2 inst_12590 ( .A(net_12004), .Z(net_12438) );
CLKBUF_X2 inst_16048 ( .A(net_15895), .Z(net_15896) );
INV_X4 inst_5581 ( .A(net_6358), .ZN(net_598) );
SDFF_X2 inst_921 ( .SI(net_8708), .Q(net_8708), .SE(net_6195), .D(net_3938), .CK(net_13020) );
CLKBUF_X2 inst_14202 ( .A(net_14049), .Z(net_14050) );
CLKBUF_X2 inst_17914 ( .A(net_17761), .Z(net_17762) );
CLKBUF_X2 inst_10772 ( .A(net_10619), .Z(net_10620) );
NAND3_X2 inst_3970 ( .A3(net_2328), .ZN(net_2251), .A1(net_2250), .A2(net_1900) );
DFFR_X1 inst_7425 ( .QN(net_8919), .D(net_4862), .CK(net_16700), .RN(x6501) );
CLKBUF_X2 inst_16633 ( .A(net_16480), .Z(net_16481) );
CLKBUF_X2 inst_11499 ( .A(net_11346), .Z(net_11347) );
INV_X2 inst_6395 ( .ZN(net_1170), .A(net_1169) );
AOI221_X2 inst_8825 ( .B1(net_8055), .C1(net_7851), .B2(net_6107), .ZN(net_6001), .C2(net_4400), .A(net_4308) );
CLKBUF_X2 inst_16273 ( .A(net_13207), .Z(net_16121) );
SDFF_X2 inst_790 ( .SI(net_8361), .Q(net_8361), .D(net_3941), .SE(net_3880), .CK(net_10332) );
CLKBUF_X2 inst_18686 ( .A(net_18533), .Z(net_18534) );
SDFF_X2 inst_1009 ( .SI(net_7311), .Q(net_6652), .D(net_6652), .SE(net_3126), .CK(net_9937) );
CLKBUF_X2 inst_10515 ( .A(net_10362), .Z(net_10363) );
AOI21_X2 inst_8931 ( .B2(net_5843), .ZN(net_5680), .A(net_5664), .B1(x338) );
AOI22_X2 inst_8024 ( .B1(net_8100), .A1(net_7760), .B2(net_6108), .A2(net_6096), .ZN(net_4113) );
CLKBUF_X2 inst_13217 ( .A(net_13064), .Z(net_13065) );
SDFF_X2 inst_733 ( .SI(net_8359), .Q(net_8359), .D(net_3954), .SE(net_3880), .CK(net_10991) );
INV_X4 inst_5885 ( .A(net_7309), .ZN(net_718) );
SDFF_X2 inst_1959 ( .D(net_7288), .SI(net_6865), .Q(net_6865), .SE(net_6282), .CK(net_14871) );
CLKBUF_X2 inst_16106 ( .A(net_15953), .Z(net_15954) );
CLKBUF_X2 inst_14294 ( .A(net_11010), .Z(net_14142) );
CLKBUF_X2 inst_16753 ( .A(net_16600), .Z(net_16601) );
AOI22_X2 inst_8020 ( .B1(net_8031), .A1(net_7997), .B2(net_6102), .A2(net_6097), .ZN(net_4116) );
AOI22_X2 inst_7892 ( .B2(net_5609), .ZN(net_4538), .A2(net_4537), .B1(net_353), .A1(net_261) );
CLKBUF_X2 inst_18162 ( .A(net_18009), .Z(net_18010) );
INV_X2 inst_6416 ( .A(net_7305), .ZN(net_839) );
CLKBUF_X2 inst_16690 ( .A(net_13801), .Z(net_16538) );
NAND2_X2 inst_4471 ( .A2(net_5463), .ZN(net_4646), .A1(net_438) );
SDFF_X2 inst_615 ( .SI(net_8378), .Q(net_8378), .D(net_3981), .SE(net_3969), .CK(net_10722) );
CLKBUF_X2 inst_12182 ( .A(net_9565), .Z(net_12030) );
CLKBUF_X2 inst_12597 ( .A(net_12444), .Z(net_12445) );
AND2_X2 inst_9157 ( .ZN(net_2833), .A1(net_2832), .A2(net_2831) );
CLKBUF_X2 inst_16877 ( .A(net_16724), .Z(net_16725) );
AOI22_X2 inst_8456 ( .B1(net_6538), .A1(net_6505), .A2(net_6137), .B2(net_6104), .ZN(net_3484) );
AOI22_X2 inst_7906 ( .B2(net_5609), .A2(net_4537), .ZN(net_4520), .A1(net_2547), .B1(net_352) );
NAND4_X2 inst_3843 ( .ZN(net_1840), .A1(net_1587), .A4(net_1559), .A2(net_1223), .A3(net_985) );
CLKBUF_X2 inst_11583 ( .A(net_10119), .Z(net_11431) );
CLKBUF_X2 inst_10621 ( .A(net_10468), .Z(net_10469) );
CLKBUF_X2 inst_17360 ( .A(net_17207), .Z(net_17208) );
CLKBUF_X2 inst_13632 ( .A(net_13479), .Z(net_13480) );
INV_X4 inst_5593 ( .A(net_6316), .ZN(net_2676) );
CLKBUF_X2 inst_10255 ( .A(net_10102), .Z(net_10103) );
MUX2_X2 inst_4941 ( .A(net_7480), .B(net_2760), .Z(net_2645), .S(net_2439) );
CLKBUF_X2 inst_18631 ( .A(net_18478), .Z(net_18479) );
AOI22_X2 inst_7835 ( .A2(net_5595), .B2(net_4881), .ZN(net_4676), .A1(net_328), .B1(net_246) );
INV_X4 inst_5133 ( .ZN(net_4353), .A(net_4315) );
DFFR_X2 inst_7095 ( .QN(net_6469), .D(net_3345), .CK(net_15111), .RN(x6501) );
CLKBUF_X2 inst_9986 ( .A(net_9833), .Z(net_9834) );
SDFFR_X2 inst_2412 ( .D(net_6320), .SE(net_2313), .SI(net_442), .Q(net_442), .CK(net_14705), .RN(x6501) );
MUX2_X2 inst_4928 ( .S(net_3537), .Z(net_3387), .B(net_3386), .A(net_602) );
CLKBUF_X2 inst_10384 ( .A(net_9528), .Z(net_10232) );
SDFFR_X2 inst_2214 ( .Q(net_7469), .D(net_7469), .SE(net_2863), .CK(net_12195), .SI(x13440), .RN(x6501) );
CLKBUF_X2 inst_18956 ( .A(net_18803), .Z(net_18804) );
CLKBUF_X2 inst_10018 ( .A(net_9523), .Z(net_9866) );
CLKBUF_X2 inst_14051 ( .A(net_13898), .Z(net_13899) );
SDFFR_X2 inst_2495 ( .Q(net_9003), .D(net_9003), .SI(net_2620), .SE(net_2562), .CK(net_16406), .RN(x6501) );
NAND2_X4 inst_4019 ( .ZN(net_4357), .A1(net_4272), .A2(net_2845) );
DFFS_X2 inst_6902 ( .QN(net_6326), .D(net_2388), .CK(net_17610), .SN(x6501) );
CLKBUF_X2 inst_11265 ( .A(net_11112), .Z(net_11113) );
CLKBUF_X2 inst_18147 ( .A(net_16530), .Z(net_17995) );
CLKBUF_X2 inst_11697 ( .A(net_9977), .Z(net_11545) );
NOR4_X2 inst_3236 ( .ZN(net_1811), .A3(net_1510), .A4(net_1418), .A2(net_1414), .A1(net_1396) );
CLKBUF_X2 inst_11219 ( .A(net_9948), .Z(net_11067) );
CLKBUF_X2 inst_10474 ( .A(net_10318), .Z(net_10322) );
CLKBUF_X2 inst_11096 ( .A(net_10490), .Z(net_10944) );
CLKBUF_X2 inst_15759 ( .A(net_15606), .Z(net_15607) );
NOR2_X2 inst_3408 ( .A2(net_6255), .A1(net_6055), .ZN(net_3574) );
XOR2_X1 inst_88 ( .Z(net_1764), .B(net_1763), .A(net_1678) );
CLKBUF_X2 inst_17369 ( .A(net_17216), .Z(net_17217) );
INV_X4 inst_6054 ( .A(net_6379), .ZN(net_495) );
CLKBUF_X2 inst_10397 ( .A(net_10244), .Z(net_10245) );
CLKBUF_X2 inst_10356 ( .A(net_9123), .Z(net_10204) );
CLKBUF_X2 inst_11190 ( .A(net_11037), .Z(net_11038) );
SDFF_X2 inst_360 ( .SI(net_8526), .Q(net_8526), .D(net_3981), .SE(net_3979), .CK(net_13011) );
CLKBUF_X2 inst_14646 ( .A(net_14493), .Z(net_14494) );
INV_X2 inst_6604 ( .A(net_6164), .ZN(net_6161) );
CLKBUF_X2 inst_10876 ( .A(net_10723), .Z(net_10724) );
CLKBUF_X2 inst_18786 ( .A(net_9419), .Z(net_18634) );
NAND3_X2 inst_3908 ( .ZN(net_5630), .A1(net_5559), .A3(net_5493), .A2(net_5362) );
CLKBUF_X2 inst_12574 ( .A(net_12421), .Z(net_12422) );
DFF_X1 inst_6797 ( .QN(net_8244), .D(net_4436), .CK(net_13591) );
SDFF_X2 inst_1129 ( .D(net_7336), .SI(net_6578), .Q(net_6578), .SE(net_3070), .CK(net_9458) );
AOI21_X2 inst_8922 ( .B2(net_5871), .ZN(net_5708), .A(net_5698), .B1(net_2727) );
SDFF_X2 inst_744 ( .Q(net_8779), .D(net_8779), .SI(net_3943), .SE(net_3879), .CK(net_13335) );
CLKBUF_X2 inst_13116 ( .A(net_10894), .Z(net_12964) );
CLKBUF_X2 inst_17104 ( .A(net_12719), .Z(net_16952) );
CLKBUF_X2 inst_13375 ( .A(net_13222), .Z(net_13223) );
NAND4_X2 inst_3827 ( .ZN(net_2747), .A2(net_2393), .A1(net_2392), .A3(x3079), .A4(x3028) );
CLKBUF_X2 inst_18720 ( .A(net_18567), .Z(net_18568) );
CLKBUF_X2 inst_12385 ( .A(net_12232), .Z(net_12233) );
CLKBUF_X2 inst_17362 ( .A(net_17209), .Z(net_17210) );
NAND2_X2 inst_4112 ( .ZN(net_5417), .A1(net_5235), .A2(net_5010) );
CLKBUF_X2 inst_13492 ( .A(net_10233), .Z(net_13340) );
CLKBUF_X2 inst_16357 ( .A(net_16204), .Z(net_16205) );
CLKBUF_X2 inst_17898 ( .A(net_17745), .Z(net_17746) );
CLKBUF_X2 inst_11002 ( .A(net_10849), .Z(net_10850) );
CLKBUF_X2 inst_15487 ( .A(net_15334), .Z(net_15335) );
SDFF_X2 inst_536 ( .Q(net_8667), .D(net_8667), .SI(net_3961), .SE(net_3935), .CK(net_13201) );
CLKBUF_X2 inst_12711 ( .A(net_12558), .Z(net_12559) );
CLKBUF_X2 inst_16243 ( .A(net_16090), .Z(net_16091) );
CLKBUF_X2 inst_11032 ( .A(net_10270), .Z(net_10880) );
SDFF_X2 inst_2027 ( .SI(net_7914), .Q(net_7914), .D(net_2708), .SE(net_2461), .CK(net_18259) );
AOI22_X2 inst_8146 ( .B1(net_8187), .A1(net_7677), .B2(net_6099), .A2(net_4399), .ZN(net_4005) );
INV_X4 inst_5882 ( .A(net_6312), .ZN(net_2667) );
DFFR_X1 inst_7487 ( .QN(net_7420), .D(net_4207), .CK(net_13382), .RN(x6501) );
SDFF_X2 inst_416 ( .SI(net_8330), .Q(net_8330), .SE(net_3978), .D(net_3976), .CK(net_12801) );
CLKBUF_X2 inst_15773 ( .A(net_15620), .Z(net_15621) );
AND2_X2 inst_9169 ( .A2(net_2553), .ZN(net_2550), .A1(net_2549) );
CLKBUF_X2 inst_10871 ( .A(net_10152), .Z(net_10719) );
SDFF_X2 inst_1406 ( .SI(net_7277), .Q(net_7134), .D(net_7134), .SE(net_6279), .CK(net_17396) );
AOI22_X2 inst_8396 ( .B1(net_8674), .A1(net_8637), .ZN(net_6236), .B2(net_6109), .A2(net_3857) );
INV_X4 inst_5500 ( .ZN(net_702), .A(x3258) );
INV_X4 inst_5330 ( .A(net_1350), .ZN(net_1349) );
NAND2_X2 inst_4319 ( .A1(net_7058), .A2(net_5162), .ZN(net_5138) );
CLKBUF_X2 inst_9520 ( .A(net_9367), .Z(net_9368) );
CLKBUF_X2 inst_10943 ( .A(net_10790), .Z(net_10791) );
CLKBUF_X2 inst_18392 ( .A(net_12986), .Z(net_18240) );
AOI22_X2 inst_8046 ( .B1(net_8137), .A1(net_7899), .A2(net_6098), .B2(net_4190), .ZN(net_4094) );
CLKBUF_X2 inst_18257 ( .A(net_18104), .Z(net_18105) );
NAND2_X2 inst_4432 ( .A1(net_6842), .A2(net_5016), .ZN(net_4995) );
CLKBUF_X2 inst_11039 ( .A(net_10886), .Z(net_10887) );
CLKBUF_X2 inst_13014 ( .A(net_12861), .Z(net_12862) );
SDFF_X2 inst_973 ( .SI(net_7336), .Q(net_6743), .D(net_6743), .SE(net_3124), .CK(net_9505) );
OAI21_X2 inst_3058 ( .B2(net_8242), .B1(net_4850), .ZN(net_4749), .A(net_2599) );
CLKBUF_X2 inst_13374 ( .A(net_13221), .Z(net_13222) );
CLKBUF_X2 inst_11258 ( .A(net_11105), .Z(net_11106) );
CLKBUF_X2 inst_11884 ( .A(net_11731), .Z(net_11732) );
CLKBUF_X2 inst_11771 ( .A(net_11618), .Z(net_11619) );
OAI21_X2 inst_3089 ( .ZN(net_2898), .B2(net_2897), .A(net_2894), .B1(net_1641) );
CLKBUF_X2 inst_18309 ( .A(net_18156), .Z(net_18157) );
SDFF_X2 inst_1122 ( .D(net_7327), .SI(net_6569), .Q(net_6569), .SE(net_3070), .CK(net_9842) );
CLKBUF_X2 inst_15009 ( .A(net_14856), .Z(net_14857) );
CLKBUF_X2 inst_12170 ( .A(net_9720), .Z(net_12018) );
NOR2_X4 inst_3324 ( .ZN(net_6079), .A2(net_5988), .A1(net_5987) );
DFFR_X1 inst_7478 ( .QN(net_7436), .D(net_4219), .CK(net_10114), .RN(x6501) );
AOI22_X2 inst_7987 ( .B1(net_8062), .A1(net_7858), .B2(net_6107), .ZN(net_6008), .A2(net_4400) );
CLKBUF_X2 inst_14351 ( .A(net_12901), .Z(net_14199) );
OAI21_X4 inst_2981 ( .B2(net_7652), .ZN(net_3301), .B1(net_3178), .A(net_3083) );
CLKBUF_X2 inst_15677 ( .A(net_15524), .Z(net_15525) );
MUX2_X2 inst_4998 ( .A(net_9038), .Z(net_3942), .B(net_3274), .S(net_622) );
CLKBUF_X2 inst_15403 ( .A(net_14304), .Z(net_15251) );
INV_X4 inst_5390 ( .ZN(net_1347), .A(net_1087) );
CLKBUF_X2 inst_9240 ( .A(net_9087), .Z(net_9088) );
NAND2_X2 inst_4406 ( .A1(net_7048), .A2(net_5162), .ZN(net_5051) );
INV_X32 inst_6169 ( .ZN(net_5164), .A(net_4815) );
HA_X1 inst_6696 ( .B(net_6105), .S(net_2820), .CO(net_2819), .A(net_2818) );
CLKBUF_X2 inst_19125 ( .A(net_18972), .Z(net_18973) );
XOR2_X1 inst_90 ( .Z(net_1665), .A(net_1567), .B(net_741) );
CLKBUF_X2 inst_11166 ( .A(net_9099), .Z(net_11014) );
CLKBUF_X2 inst_14950 ( .A(net_14797), .Z(net_14798) );
CLKBUF_X2 inst_16348 ( .A(net_11389), .Z(net_16196) );
CLKBUF_X2 inst_17875 ( .A(net_17722), .Z(net_17723) );
DFF_X1 inst_6858 ( .Q(net_6445), .D(net_3623), .CK(net_17888) );
CLKBUF_X2 inst_10850 ( .A(net_10697), .Z(net_10698) );
CLKBUF_X2 inst_18910 ( .A(net_18757), .Z(net_18758) );
NAND2_X2 inst_4650 ( .ZN(net_2467), .A1(net_2307), .A2(net_2153) );
AOI221_X2 inst_8860 ( .ZN(net_2249), .A(net_2248), .C1(net_2247), .C2(net_2172), .B1(net_1283), .B2(net_1063) );
DFFR_X2 inst_7197 ( .D(net_2363), .QN(net_212), .CK(net_15011), .RN(x6501) );
INV_X4 inst_5093 ( .ZN(net_5704), .A(net_5680) );
NAND4_X2 inst_3833 ( .ZN(net_2291), .A4(net_2018), .A3(net_1811), .A1(net_1406), .A2(net_1392) );
SDFFR_X2 inst_2460 ( .SE(net_2748), .D(net_2640), .SI(net_456), .Q(net_456), .CK(net_13926), .RN(x6501) );
AOI22_X2 inst_8457 ( .B1(net_6737), .A1(net_6704), .B2(net_6202), .A2(net_3520), .ZN(net_3483) );
CLKBUF_X2 inst_18893 ( .A(net_18740), .Z(net_18741) );
SDFF_X2 inst_1217 ( .Q(net_7815), .D(net_7815), .SE(net_2730), .SI(net_2573), .CK(net_18098) );
CLKBUF_X2 inst_15936 ( .A(net_15783), .Z(net_15784) );
CLKBUF_X2 inst_10832 ( .A(net_10679), .Z(net_10680) );
CLKBUF_X2 inst_18706 ( .A(net_18553), .Z(net_18554) );
CLKBUF_X2 inst_10788 ( .A(net_10158), .Z(net_10636) );
CLKBUF_X2 inst_16372 ( .A(net_16219), .Z(net_16220) );
CLKBUF_X2 inst_10285 ( .A(net_10132), .Z(net_10133) );
DFFS_X1 inst_6938 ( .D(net_6145), .CK(net_13650), .SN(x6501), .Q(x725) );
DFFR_X2 inst_7126 ( .Q(net_7353), .D(net_3066), .CK(net_9650), .RN(x6501) );
CLKBUF_X2 inst_10187 ( .A(net_10034), .Z(net_10035) );
CLKBUF_X2 inst_15545 ( .A(net_15392), .Z(net_15393) );
OAI21_X2 inst_3027 ( .B2(net_8234), .B1(net_4954), .ZN(net_4944), .A(net_4832) );
INV_X4 inst_5907 ( .ZN(net_2701), .A(net_267) );
CLKBUF_X2 inst_17762 ( .A(net_17609), .Z(net_17610) );
AOI222_X1 inst_8614 ( .B2(net_6760), .B1(net_5835), .A2(net_5830), .C2(net_5824), .ZN(net_5799), .C1(net_2145), .A1(net_1675) );
CLKBUF_X2 inst_14016 ( .A(net_11484), .Z(net_13864) );
CLKBUF_X2 inst_14059 ( .A(net_13906), .Z(net_13907) );
CLKBUF_X2 inst_18283 ( .A(net_12649), .Z(net_18131) );
CLKBUF_X2 inst_10235 ( .A(net_10082), .Z(net_10083) );
CLKBUF_X2 inst_15843 ( .A(net_15690), .Z(net_15691) );
DFFR_X1 inst_7480 ( .QN(net_7423), .D(net_4212), .CK(net_12316), .RN(x6501) );
XOR2_X1 inst_68 ( .Z(net_3991), .B(net_3990), .A(net_3582) );
AOI22_X2 inst_8029 ( .B1(net_8169), .A1(net_7727), .B2(net_6101), .A2(net_6095), .ZN(net_6018) );
CLKBUF_X2 inst_18725 ( .A(net_18572), .Z(net_18573) );
CLKBUF_X2 inst_18289 ( .A(net_18136), .Z(net_18137) );
SDFF_X2 inst_1253 ( .SI(net_7674), .Q(net_7674), .SE(net_2714), .D(net_2709), .CK(net_18583) );
CLKBUF_X2 inst_10913 ( .A(net_9826), .Z(net_10761) );
CLKBUF_X2 inst_10689 ( .A(net_10536), .Z(net_10537) );
CLKBUF_X2 inst_11943 ( .A(net_11790), .Z(net_11791) );
OR4_X2 inst_2793 ( .A4(net_3542), .ZN(net_2458), .A1(net_2306), .A2(net_534), .A3(x3762) );
CLKBUF_X2 inst_15647 ( .A(net_9972), .Z(net_15495) );
SDFF_X2 inst_2018 ( .SI(net_7774), .Q(net_7774), .D(net_2705), .SE(net_2459), .CK(net_18509) );
SDFF_X2 inst_1884 ( .D(net_7295), .SI(net_6992), .Q(net_6992), .SE(net_6283), .CK(net_15407) );
INV_X2 inst_6488 ( .A(net_7574), .ZN(net_3142) );
CLKBUF_X2 inst_13172 ( .A(net_13019), .Z(net_13020) );
AOI22_X2 inst_8540 ( .B1(net_6527), .A1(net_6494), .A2(net_6137), .B2(net_6104), .ZN(net_3400) );
SDFF_X2 inst_1690 ( .Q(net_8020), .D(net_8020), .SI(net_2584), .SE(net_2545), .CK(net_16030) );
INV_X2 inst_6413 ( .ZN(net_870), .A(net_869) );
CLKBUF_X2 inst_9815 ( .A(net_9662), .Z(net_9663) );
INV_X4 inst_5312 ( .ZN(net_2043), .A(net_1136) );
CLKBUF_X2 inst_9540 ( .A(net_9344), .Z(net_9388) );
CLKBUF_X2 inst_13015 ( .A(net_12862), .Z(net_12863) );
SDFF_X2 inst_1287 ( .Q(net_8107), .D(net_8107), .SE(net_2707), .SI(net_2660), .CK(net_17093) );
NAND2_X2 inst_4231 ( .A1(net_6899), .A2(net_5247), .ZN(net_5229) );
CLKBUF_X2 inst_16840 ( .A(net_16687), .Z(net_16688) );
CLKBUF_X2 inst_17333 ( .A(net_17180), .Z(net_17181) );
SDFF_X2 inst_1169 ( .D(net_7335), .SI(net_6511), .Q(net_6511), .SE(net_3071), .CK(net_9747) );
NAND2_X2 inst_4266 ( .A1(net_7035), .A2(net_5249), .ZN(net_5194) );
INV_X4 inst_5826 ( .A(net_7422), .ZN(net_2818) );
NOR2_X2 inst_3483 ( .ZN(net_2235), .A1(net_2234), .A2(net_2233) );
CLKBUF_X2 inst_17921 ( .A(net_17768), .Z(net_17769) );
INV_X4 inst_5704 ( .A(net_7254), .ZN(net_1958) );
AOI222_X1 inst_8634 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_4276), .B1(net_3922), .C1(net_3921), .A1(x13633) );
CLKBUF_X2 inst_9440 ( .A(net_9264), .Z(net_9288) );
CLKBUF_X2 inst_17522 ( .A(net_17369), .Z(net_17370) );
CLKBUF_X2 inst_12251 ( .A(net_12098), .Z(net_12099) );
CLKBUF_X2 inst_17788 ( .A(net_17635), .Z(net_17636) );
OR2_X2 inst_2877 ( .ZN(net_3530), .A2(net_3529), .A1(net_3526) );
CLKBUF_X2 inst_12908 ( .A(net_12755), .Z(net_12756) );
CLKBUF_X2 inst_15150 ( .A(net_12058), .Z(net_14998) );
CLKBUF_X2 inst_16331 ( .A(net_16178), .Z(net_16179) );
INV_X2 inst_6514 ( .A(net_8950), .ZN(net_753) );
CLKBUF_X2 inst_11221 ( .A(net_9729), .Z(net_11069) );
CLKBUF_X2 inst_16561 ( .A(net_16408), .Z(net_16409) );
DFFR_X1 inst_7502 ( .QN(net_6336), .D(net_1896), .CK(net_17800), .RN(x6501) );
CLKBUF_X2 inst_11709 ( .A(net_11556), .Z(net_11557) );
CLKBUF_X2 inst_12062 ( .A(net_11909), .Z(net_11910) );
CLKBUF_X2 inst_18983 ( .A(net_15742), .Z(net_18831) );
SDFF_X2 inst_1418 ( .SI(net_7297), .Q(net_7074), .D(net_7074), .SE(net_6280), .CK(net_15457) );
AND2_X4 inst_9095 ( .ZN(net_2538), .A1(net_2274), .A2(net_2268) );
CLKBUF_X2 inst_14124 ( .A(net_13849), .Z(net_13972) );
SDFF_X2 inst_1740 ( .Q(net_7878), .D(net_7878), .SI(net_2709), .SE(net_2543), .CK(net_15741) );
CLKBUF_X2 inst_10171 ( .A(net_9750), .Z(net_10019) );
CLKBUF_X2 inst_14499 ( .A(net_14346), .Z(net_14347) );
INV_X4 inst_5663 ( .A(net_7389), .ZN(net_1033) );
CLKBUF_X2 inst_16126 ( .A(net_15973), .Z(net_15974) );
CLKBUF_X2 inst_16433 ( .A(net_14689), .Z(net_16281) );
AOI22_X2 inst_7822 ( .B1(net_7513), .A2(net_5535), .B2(net_5260), .ZN(net_4702), .A1(net_472) );
CLKBUF_X2 inst_11176 ( .A(net_10609), .Z(net_11024) );
SDFF_X2 inst_2001 ( .SI(net_7789), .Q(net_7789), .D(net_2719), .SE(net_2459), .CK(net_18739) );
NAND2_X2 inst_4836 ( .ZN(net_988), .A1(net_613), .A2(net_612) );
CLKBUF_X2 inst_18602 ( .A(net_18449), .Z(net_18450) );
SDFF_X2 inst_1657 ( .SI(net_7738), .Q(net_7738), .D(net_2721), .SE(net_2560), .CK(net_15753) );
CLKBUF_X2 inst_10321 ( .A(net_10168), .Z(net_10169) );
CLKBUF_X2 inst_12982 ( .A(net_12829), .Z(net_12830) );
CLKBUF_X2 inst_14385 ( .A(net_14232), .Z(net_14233) );
CLKBUF_X2 inst_15570 ( .A(net_15417), .Z(net_15418) );
SDFFS_X2 inst_2077 ( .SI(net_7382), .SE(net_2795), .Q(net_171), .D(net_171), .CK(net_17497), .SN(x6501) );
CLKBUF_X2 inst_10085 ( .A(net_9932), .Z(net_9933) );
CLKBUF_X2 inst_17057 ( .A(net_16904), .Z(net_16905) );
CLKBUF_X2 inst_14473 ( .A(net_14320), .Z(net_14321) );
AOI22_X2 inst_8078 ( .B1(net_8012), .A1(net_7978), .B2(net_6102), .A2(net_6097), .ZN(net_6048) );
CLKBUF_X2 inst_12729 ( .A(net_10028), .Z(net_12577) );
CLKBUF_X2 inst_13704 ( .A(net_12551), .Z(net_13552) );
CLKBUF_X2 inst_13930 ( .A(net_13777), .Z(net_13778) );
INV_X1 inst_6656 ( .A(net_6169), .ZN(net_6167) );
CLKBUF_X2 inst_12179 ( .A(net_9309), .Z(net_12027) );
SDFF_X2 inst_1495 ( .SI(net_7851), .Q(net_7851), .D(net_2706), .SE(net_2558), .CK(net_15289) );
SDFF_X2 inst_797 ( .SI(net_8369), .Q(net_8369), .D(net_3949), .SE(net_3880), .CK(net_12584) );
INV_X8 inst_5051 ( .ZN(net_6194), .A(net_6190) );
INV_X4 inst_5546 ( .A(net_1809), .ZN(net_641) );
CLKBUF_X2 inst_9310 ( .A(net_9157), .Z(net_9158) );
CLKBUF_X2 inst_17318 ( .A(net_17165), .Z(net_17166) );
OAI21_X2 inst_3032 ( .ZN(net_4854), .B2(net_4853), .B1(net_4850), .A(net_2623) );
AOI21_X2 inst_8882 ( .ZN(net_5922), .A(net_5783), .B2(net_5749), .B1(net_4903) );
CLKBUF_X2 inst_17489 ( .A(net_17336), .Z(net_17337) );
CLKBUF_X2 inst_12069 ( .A(net_11916), .Z(net_11917) );
DFF_X1 inst_6856 ( .QN(net_6444), .D(net_3625), .CK(net_17889) );
DFF_X1 inst_6787 ( .Q(net_7536), .D(net_4583), .CK(net_11953) );
CLKBUF_X2 inst_13195 ( .A(net_13042), .Z(net_13043) );
CLKBUF_X2 inst_14699 ( .A(net_13675), .Z(net_14547) );
NOR2_X2 inst_3583 ( .ZN(net_3320), .A1(net_1075), .A2(net_1074) );
CLKBUF_X2 inst_13242 ( .A(net_12460), .Z(net_13090) );
AOI22_X2 inst_8446 ( .B1(net_6668), .A1(net_6635), .A2(net_6213), .B2(net_6138), .ZN(net_3494) );
SDFF_X2 inst_1115 ( .D(net_7318), .SI(net_6527), .Q(net_6527), .SE(net_3086), .CK(net_9917) );
MUX2_X2 inst_4933 ( .B(net_8894), .S(net_3153), .Z(net_3034), .A(net_1459) );
CLKBUF_X2 inst_17793 ( .A(net_12686), .Z(net_17641) );
INV_X2 inst_6234 ( .ZN(net_5476), .A(net_5290) );
SDFF_X2 inst_1021 ( .SI(net_7337), .Q(net_6678), .D(net_6678), .SE(net_3126), .CK(net_9492) );
OAI221_X2 inst_2976 ( .C2(net_7169), .B2(net_7168), .ZN(net_2028), .B1(net_1830), .C1(net_1829), .A(net_1652) );
CLKBUF_X2 inst_17662 ( .A(net_17509), .Z(net_17510) );
AND2_X4 inst_9140 ( .ZN(net_1381), .A2(net_787), .A1(net_176) );
NAND2_X2 inst_4204 ( .ZN(net_5292), .A2(net_5174), .A1(net_5051) );
CLKBUF_X2 inst_18116 ( .A(net_17963), .Z(net_17964) );
CLKBUF_X2 inst_12095 ( .A(net_11942), .Z(net_11943) );
NAND2_X2 inst_4827 ( .A2(net_7305), .ZN(net_1352), .A1(net_655) );
SDFF_X2 inst_572 ( .Q(net_8836), .D(net_8836), .SE(net_3964), .SI(net_3956), .CK(net_10065) );
CLKBUF_X2 inst_12699 ( .A(net_11686), .Z(net_12547) );
CLKBUF_X2 inst_12392 ( .A(net_12239), .Z(net_12240) );
XNOR2_X2 inst_257 ( .B(net_2684), .A(net_2682), .ZN(net_1190) );
INV_X8 inst_5036 ( .ZN(net_6092), .A(net_3575) );
CLKBUF_X2 inst_15062 ( .A(net_9898), .Z(net_14910) );
CLKBUF_X2 inst_17449 ( .A(net_13026), .Z(net_17297) );
SDFF_X2 inst_485 ( .SI(net_8608), .Q(net_8608), .SE(net_3984), .D(net_3973), .CK(net_13205) );
CLKBUF_X2 inst_12971 ( .A(net_9805), .Z(net_12819) );
CLKBUF_X2 inst_10684 ( .A(net_10187), .Z(net_10532) );
CLKBUF_X2 inst_14655 ( .A(net_9339), .Z(net_14503) );
SDFF_X2 inst_1205 ( .Q(net_7974), .D(net_7974), .SE(net_2755), .SI(net_2656), .CK(net_16887) );
CLKBUF_X2 inst_17609 ( .A(net_17456), .Z(net_17457) );
CLKBUF_X2 inst_18043 ( .A(net_16705), .Z(net_17891) );
INV_X4 inst_5085 ( .ZN(net_5729), .A(net_5708) );
CLKBUF_X2 inst_16286 ( .A(net_11288), .Z(net_16134) );
CLKBUF_X2 inst_11048 ( .A(net_10895), .Z(net_10896) );
CLKBUF_X2 inst_18558 ( .A(net_18405), .Z(net_18406) );
CLKBUF_X2 inst_17064 ( .A(net_16911), .Z(net_16912) );
AOI22_X2 inst_8310 ( .B1(net_8696), .A1(net_8659), .B2(net_6109), .A2(net_3857), .ZN(net_3735) );
CLKBUF_X2 inst_15012 ( .A(net_14859), .Z(net_14860) );
AOI222_X1 inst_8641 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3932), .B1(net_3229), .C1(net_3227), .A1(x13705) );
CLKBUF_X2 inst_14409 ( .A(net_14256), .Z(net_14257) );
DFFS_X1 inst_6929 ( .D(net_6145), .CK(net_16361), .SN(x6501), .Q(x852) );
NAND4_X2 inst_3716 ( .A4(net_6234), .A1(net_6233), .ZN(net_4421), .A2(net_3659), .A3(net_3658) );
CLKBUF_X2 inst_15903 ( .A(net_15750), .Z(net_15751) );
XNOR2_X2 inst_253 ( .A(net_2690), .B(net_2640), .ZN(net_1196) );
CLKBUF_X2 inst_16239 ( .A(net_14816), .Z(net_16087) );
CLKBUF_X2 inst_16219 ( .A(net_16066), .Z(net_16067) );
CLKBUF_X2 inst_14080 ( .A(net_13927), .Z(net_13928) );
CLKBUF_X2 inst_16052 ( .A(net_15899), .Z(net_15900) );
SDFF_X2 inst_589 ( .SI(net_8371), .Q(net_8371), .SE(net_3969), .D(net_3961), .CK(net_10012) );
INV_X4 inst_5229 ( .ZN(net_5522), .A(net_2252) );
CLKBUF_X2 inst_18671 ( .A(net_18518), .Z(net_18519) );
NAND2_X2 inst_4868 ( .A2(net_7405), .ZN(net_1431), .A1(net_716) );
CLKBUF_X2 inst_10176 ( .A(net_10023), .Z(net_10024) );
CLKBUF_X2 inst_11969 ( .A(net_9266), .Z(net_11817) );
NAND2_X2 inst_4273 ( .A1(net_6918), .A2(net_5247), .ZN(net_5187) );
CLKBUF_X2 inst_18461 ( .A(net_18308), .Z(net_18309) );
CLKBUF_X2 inst_17347 ( .A(net_17194), .Z(net_17195) );
CLKBUF_X2 inst_9829 ( .A(net_9676), .Z(net_9677) );
CLKBUF_X2 inst_9822 ( .A(net_9669), .Z(net_9670) );
SDFF_X2 inst_1877 ( .D(net_7284), .SI(net_6981), .Q(net_6981), .SE(net_6283), .CK(net_16187) );
XOR2_X2 inst_59 ( .A(net_3167), .Z(net_954), .B(net_581) );
SDFFR_X2 inst_2367 ( .SE(net_2260), .Q(net_323), .D(net_323), .CK(net_10463), .RN(x6501), .SI(x2981) );
AND2_X2 inst_9182 ( .ZN(net_2009), .A1(net_2008), .A2(net_2007) );
CLKBUF_X2 inst_10533 ( .A(net_10380), .Z(net_10381) );
NOR3_X2 inst_3256 ( .ZN(net_5020), .A3(net_4956), .A1(net_4927), .A2(net_3262) );
AND3_X2 inst_9050 ( .A1(net_2666), .A2(net_2569), .ZN(net_1265), .A3(net_816) );
CLKBUF_X2 inst_12867 ( .A(net_12714), .Z(net_12715) );
SDFF_X2 inst_1865 ( .D(net_7290), .SI(net_6907), .Q(net_6907), .SE(net_6284), .CK(net_15327) );
CLKBUF_X2 inst_15715 ( .A(net_15562), .Z(net_15563) );
XOR2_X2 inst_37 ( .Z(net_1119), .A(net_1118), .B(net_1117) );
INV_X2 inst_6390 ( .A(net_1925), .ZN(net_1535) );
CLKBUF_X2 inst_11960 ( .A(net_11807), .Z(net_11808) );
SDFF_X2 inst_1664 ( .SI(net_7758), .Q(net_7758), .D(net_2718), .SE(net_2560), .CK(net_18769) );
SDFF_X2 inst_1447 ( .SI(net_7296), .Q(net_7113), .D(net_7113), .SE(net_6278), .CK(net_15454) );
CLKBUF_X2 inst_14881 ( .A(net_11282), .Z(net_14729) );
CLKBUF_X2 inst_9601 ( .A(net_9059), .Z(net_9449) );
NAND2_X2 inst_4730 ( .ZN(net_2709), .A2(net_1586), .A1(net_1122) );
OAI21_X2 inst_3075 ( .B1(net_7632), .ZN(net_3903), .A(net_3902), .B2(net_3901) );
OR3_X4 inst_2800 ( .A3(net_3535), .ZN(net_3354), .A1(net_2306), .A2(x3762) );
CLKBUF_X2 inst_9487 ( .A(net_9162), .Z(net_9335) );
SDFF_X2 inst_766 ( .Q(net_8809), .D(net_8809), .SI(net_3951), .SE(net_3879), .CK(net_10594) );
SDFF_X2 inst_1908 ( .D(net_7269), .SI(net_6846), .Q(net_6846), .SE(net_6282), .CK(net_14084) );
NOR3_X2 inst_3270 ( .ZN(net_2417), .A1(net_2400), .A2(net_2397), .A3(net_2396) );
CLKBUF_X2 inst_14879 ( .A(net_14726), .Z(net_14727) );
CLKBUF_X2 inst_15957 ( .A(net_15804), .Z(net_15805) );
NOR3_X2 inst_3273 ( .A1(net_2415), .ZN(net_2413), .A3(net_2397), .A2(net_1779) );
INV_X4 inst_6139 ( .A(net_6118), .ZN(net_6116) );
CLKBUF_X2 inst_9943 ( .A(net_9790), .Z(net_9791) );
CLKBUF_X2 inst_14282 ( .A(net_14129), .Z(net_14130) );
INV_X2 inst_6552 ( .A(net_7583), .ZN(net_3137) );
SDFF_X2 inst_1619 ( .Q(net_8161), .D(net_8161), .SI(net_2576), .SE(net_2538), .CK(net_16041) );
CLKBUF_X2 inst_15344 ( .A(net_15191), .Z(net_15192) );
SDFF_X2 inst_441 ( .Q(net_8770), .D(net_8770), .SE(net_3982), .SI(net_3952), .CK(net_10378) );
OAI21_X2 inst_3110 ( .B1(net_2698), .A(net_2480), .B2(net_2479), .ZN(net_2478) );
CLKBUF_X2 inst_19001 ( .A(net_18848), .Z(net_18849) );
INV_X2 inst_6201 ( .ZN(net_5509), .A(net_5425) );
AOI22_X2 inst_8425 ( .B1(net_6729), .A1(net_6696), .B2(net_6202), .A2(net_3520), .ZN(net_3516) );
CLKBUF_X2 inst_11414 ( .A(net_10581), .Z(net_11262) );
INV_X4 inst_5228 ( .ZN(net_5783), .A(net_2252) );
CLKBUF_X2 inst_16256 ( .A(net_10657), .Z(net_16104) );
SDFF_X2 inst_808 ( .SI(net_8497), .Q(net_8497), .D(net_3973), .SE(net_3884), .CK(net_13170) );
CLKBUF_X2 inst_18622 ( .A(net_15016), .Z(net_18470) );
NAND4_X2 inst_3859 ( .A1(net_2832), .A4(net_2754), .A3(net_2494), .ZN(net_2457), .A2(net_1055) );
CLKBUF_X2 inst_18159 ( .A(net_18006), .Z(net_18007) );
CLKBUF_X2 inst_9683 ( .A(net_9530), .Z(net_9531) );
CLKBUF_X2 inst_16068 ( .A(net_15915), .Z(net_15916) );
SDFF_X2 inst_1383 ( .SI(net_7270), .Q(net_7087), .D(net_7087), .SE(net_6278), .CK(net_16868) );
OR2_X4 inst_2838 ( .ZN(net_2288), .A1(net_2287), .A2(net_2223) );
INV_X4 inst_6153 ( .A(net_6183), .ZN(net_6181) );
OR2_X4 inst_2833 ( .A2(net_6199), .A1(net_6106), .ZN(net_5902) );
NOR2_X2 inst_3423 ( .ZN(net_3095), .A2(net_3093), .A1(net_2812) );
CLKBUF_X2 inst_15349 ( .A(net_15196), .Z(net_15197) );
CLKBUF_X2 inst_16212 ( .A(net_16059), .Z(net_16060) );
SDFF_X2 inst_2042 ( .SI(net_7773), .Q(net_7773), .D(net_2585), .SE(net_2459), .CK(net_15724) );
AOI22_X2 inst_8383 ( .A1(net_8598), .B1(net_8413), .A2(net_3864), .B2(net_3863), .ZN(net_3665) );
CLKBUF_X2 inst_16070 ( .A(net_15917), .Z(net_15918) );
AOI22_X2 inst_8248 ( .B1(net_8835), .A1(net_8354), .A2(net_6265), .B2(net_6253), .ZN(net_3788) );
CLKBUF_X2 inst_19186 ( .A(net_19033), .Z(net_19034) );
CLKBUF_X2 inst_15503 ( .A(net_12738), .Z(net_15351) );
INV_X4 inst_5156 ( .ZN(net_3175), .A(net_3152) );
CLKBUF_X2 inst_13361 ( .A(net_13208), .Z(net_13209) );
CLKBUF_X2 inst_15383 ( .A(net_9934), .Z(net_15231) );
INV_X4 inst_6107 ( .A(net_7206), .ZN(net_632) );
CLKBUF_X2 inst_10758 ( .A(net_10605), .Z(net_10606) );
OR3_X4 inst_2796 ( .A1(net_4406), .ZN(net_4381), .A2(net_4380), .A3(net_4316) );
SDFFR_X1 inst_2729 ( .SI(net_9042), .Q(net_9042), .D(net_7471), .SE(net_3208), .CK(net_12216), .RN(x6501) );
CLKBUF_X2 inst_10587 ( .A(net_9287), .Z(net_10435) );
AOI22_X2 inst_8364 ( .B1(net_8814), .A1(net_8555), .A2(net_3861), .B2(net_3860), .ZN(net_3684) );
AOI221_X2 inst_8842 ( .B1(net_8050), .C1(net_7846), .B2(net_6107), .ZN(net_6029), .C2(net_4400), .A(net_4280) );
SDFF_X2 inst_1815 ( .D(net_7296), .SI(net_6953), .Q(net_6953), .SE(net_6281), .CK(net_15812) );
INV_X4 inst_5267 ( .A(net_2401), .ZN(net_1715) );
CLKBUF_X2 inst_13187 ( .A(net_13034), .Z(net_13035) );
CLKBUF_X2 inst_10422 ( .A(net_10269), .Z(net_10270) );
CLKBUF_X2 inst_16826 ( .A(net_16673), .Z(net_16674) );
CLKBUF_X2 inst_16788 ( .A(net_16635), .Z(net_16636) );
DFFR_X2 inst_7010 ( .QN(net_6295), .D(net_5754), .CK(net_16751), .RN(x6501) );
CLKBUF_X2 inst_17850 ( .A(net_17697), .Z(net_17698) );
CLKBUF_X2 inst_12379 ( .A(net_10818), .Z(net_12227) );
HA_X1 inst_6708 ( .A(net_8945), .S(net_1488), .CO(net_1487), .B(net_1274) );
CLKBUF_X2 inst_10840 ( .A(net_10687), .Z(net_10688) );
CLKBUF_X2 inst_10319 ( .A(net_9236), .Z(net_10167) );
INV_X4 inst_5442 ( .ZN(net_1134), .A(net_820) );
CLKBUF_X2 inst_17555 ( .A(net_13955), .Z(net_17403) );
NAND2_X2 inst_4758 ( .ZN(net_1737), .A2(net_1736), .A1(net_842) );
CLKBUF_X2 inst_9857 ( .A(net_9149), .Z(net_9705) );
NAND3_X4 inst_3875 ( .A1(net_6168), .A2(net_3535), .ZN(net_2210), .A3(net_2027) );
CLKBUF_X2 inst_15187 ( .A(net_15034), .Z(net_15035) );
SDFFR_X2 inst_2629 ( .Q(net_7384), .D(net_7384), .SE(net_1136), .CK(net_14952), .RN(x6501), .SI(x4667) );
AOI21_X2 inst_8989 ( .ZN(net_1707), .B2(net_1482), .B1(net_1348), .A(net_1327) );
CLKBUF_X2 inst_16421 ( .A(net_16268), .Z(net_16269) );
CLKBUF_X2 inst_13658 ( .A(net_13505), .Z(net_13506) );
CLKBUF_X2 inst_9732 ( .A(net_9579), .Z(net_9580) );
CLKBUF_X2 inst_14342 ( .A(net_9801), .Z(net_14190) );
CLKBUF_X2 inst_9595 ( .A(net_9442), .Z(net_9443) );
DFFR_X2 inst_7235 ( .QN(net_7207), .D(net_2174), .CK(net_17999), .RN(x6501) );
SDFF_X2 inst_1341 ( .Q(net_7895), .D(net_7895), .SI(net_2713), .SE(net_2543), .CK(net_14432) );
SDFF_X2 inst_587 ( .Q(net_8823), .D(net_8823), .SE(net_3964), .SI(net_3937), .CK(net_10729) );
SDFF_X2 inst_666 ( .Q(net_8441), .D(net_8441), .SI(net_3976), .SE(net_3934), .CK(net_10352) );
CLKBUF_X2 inst_10798 ( .A(net_10645), .Z(net_10646) );
CLKBUF_X2 inst_18673 ( .A(net_18520), .Z(net_18521) );
INV_X4 inst_5937 ( .A(net_6400), .ZN(net_2551) );
DFFR_X2 inst_7182 ( .QN(net_8957), .D(net_2484), .CK(net_15077), .RN(x6501) );
SDFF_X2 inst_1829 ( .D(net_7289), .SI(net_6866), .Q(net_6866), .SE(net_6282), .CK(net_15335) );
INV_X2 inst_6446 ( .ZN(net_600), .A(net_389) );
CLKBUF_X2 inst_9868 ( .A(net_9715), .Z(net_9716) );
DFFR_X1 inst_7368 ( .D(net_5937), .CK(net_11985), .RN(x6501), .Q(x1039) );
CLKBUF_X2 inst_12376 ( .A(net_12223), .Z(net_12224) );
INV_X4 inst_5252 ( .A(net_2073), .ZN(net_1833) );
CLKBUF_X2 inst_11217 ( .A(net_11064), .Z(net_11065) );
CLKBUF_X2 inst_11939 ( .A(net_11786), .Z(net_11787) );
CLKBUF_X2 inst_12210 ( .A(net_12057), .Z(net_12058) );
CLKBUF_X2 inst_13547 ( .A(net_13394), .Z(net_13395) );
CLKBUF_X2 inst_19052 ( .A(net_16691), .Z(net_18900) );
CLKBUF_X2 inst_17507 ( .A(net_17354), .Z(net_17355) );
NOR3_X2 inst_3315 ( .ZN(net_2156), .A3(net_1430), .A1(net_1178), .A2(net_914) );
DFFR_X2 inst_7347 ( .Q(net_7323), .CK(net_11770), .D(x13069), .RN(x6501) );
AOI22_X2 inst_7753 ( .B1(net_6981), .A1(net_6941), .A2(net_5443), .B2(net_5442), .ZN(net_5394) );
CLKBUF_X2 inst_15783 ( .A(net_15630), .Z(net_15631) );
CLKBUF_X2 inst_18426 ( .A(net_18092), .Z(net_18274) );
CLKBUF_X2 inst_11652 ( .A(net_10247), .Z(net_11500) );
CLKBUF_X2 inst_13094 ( .A(net_10949), .Z(net_12942) );
CLKBUF_X2 inst_14809 ( .A(net_14656), .Z(net_14657) );
SDFF_X2 inst_343 ( .SI(net_8451), .Q(net_8451), .SE(net_3983), .D(net_3947), .CK(net_12485) );
CLKBUF_X2 inst_10431 ( .A(net_10278), .Z(net_10279) );
NAND2_X2 inst_4739 ( .ZN(net_2590), .A2(net_1586), .A1(net_945) );
SDFF_X2 inst_1106 ( .D(net_7337), .SI(net_6546), .Q(net_6546), .SE(net_3086), .CK(net_9468) );
SDFF_X2 inst_543 ( .Q(net_8668), .D(net_8668), .SI(net_3943), .SE(net_3935), .CK(net_13351) );
CLKBUF_X2 inst_12131 ( .A(net_11978), .Z(net_11979) );
CLKBUF_X2 inst_14194 ( .A(net_14041), .Z(net_14042) );
DFFS_X2 inst_6882 ( .Q(net_8261), .D(net_3120), .CK(net_18476), .SN(x6501) );
CLKBUF_X2 inst_13122 ( .A(net_9643), .Z(net_12970) );
CLKBUF_X2 inst_16915 ( .A(net_16762), .Z(net_16763) );
SDFFS_X2 inst_2070 ( .SI(net_7379), .SE(net_2794), .Q(net_168), .D(net_168), .CK(net_17740), .SN(x6501) );
OR2_X2 inst_2890 ( .A1(net_2263), .A2(net_2261), .ZN(net_1579) );
INV_X4 inst_5765 ( .A(net_7480), .ZN(net_1656) );
CLKBUF_X2 inst_13858 ( .A(net_13705), .Z(net_13706) );
INV_X2 inst_6337 ( .ZN(net_2857), .A(net_2792) );
CLKBUF_X2 inst_12538 ( .A(net_11705), .Z(net_12386) );
CLKBUF_X2 inst_18292 ( .A(net_18139), .Z(net_18140) );
CLKBUF_X2 inst_16109 ( .A(net_15956), .Z(net_15957) );
DFFR_X1 inst_7555 ( .Q(net_8288), .D(net_8278), .CK(net_12229), .RN(x6501) );
AOI22_X2 inst_8347 ( .B1(net_8701), .A1(net_8664), .ZN(net_6238), .B2(net_6109), .A2(net_3857) );
NAND2_X2 inst_4304 ( .A1(net_7053), .A2(net_5162), .ZN(net_5153) );
DFF_X1 inst_6848 ( .Q(net_6436), .D(net_3633), .CK(net_17906) );
SDFFR_X1 inst_2745 ( .SI(net_9044), .Q(net_9044), .D(net_7473), .SE(net_3208), .CK(net_12204), .RN(x6501) );
CLKBUF_X2 inst_13810 ( .A(net_9663), .Z(net_13658) );
CLKBUF_X2 inst_16719 ( .A(net_16566), .Z(net_16567) );
DFFR_X2 inst_7253 ( .QN(net_7227), .D(net_2062), .CK(net_15042), .RN(x6501) );
CLKBUF_X2 inst_11802 ( .A(net_11649), .Z(net_11650) );
CLKBUF_X2 inst_11297 ( .A(net_11144), .Z(net_11145) );
CLKBUF_X2 inst_13125 ( .A(net_12972), .Z(net_12973) );
CLKBUF_X2 inst_12452 ( .A(net_12299), .Z(net_12300) );
CLKBUF_X2 inst_15959 ( .A(net_15806), .Z(net_15807) );
SDFF_X2 inst_1244 ( .SI(net_7670), .Q(net_7670), .D(net_2721), .SE(net_2714), .CK(net_18588) );
NAND2_X2 inst_4410 ( .A1(net_6840), .ZN(net_5018), .A2(net_5016) );
AOI22_X2 inst_8134 ( .B1(net_8084), .A1(net_7744), .B2(net_6108), .A2(net_6096), .ZN(net_4016) );
SDFF_X2 inst_582 ( .Q(net_8849), .D(net_8849), .SE(net_3964), .SI(net_3939), .CK(net_10551) );
NAND2_X2 inst_4515 ( .ZN(net_4227), .A1(net_3881), .A2(net_3337) );
SDFF_X2 inst_1850 ( .D(net_7272), .SI(net_6889), .Q(net_6889), .SE(net_6284), .CK(net_14110) );
NOR2_X2 inst_3477 ( .A1(net_3023), .ZN(net_2301), .A2(net_2228) );
SDFF_X2 inst_1950 ( .D(net_7276), .SI(net_6933), .Q(net_6933), .SE(net_6281), .CK(net_17340) );
CLKBUF_X2 inst_12057 ( .A(net_11904), .Z(net_11905) );
INV_X4 inst_5287 ( .ZN(net_1784), .A(net_1379) );
CLKBUF_X2 inst_9402 ( .A(net_9249), .Z(net_9250) );
CLKBUF_X2 inst_16606 ( .A(net_16453), .Z(net_16454) );
DFFR_X2 inst_7292 ( .D(net_399), .QN(net_396), .CK(net_18716), .RN(x6501) );
CLKBUF_X2 inst_12673 ( .A(net_10012), .Z(net_12521) );
CLKBUF_X2 inst_14727 ( .A(net_9969), .Z(net_14575) );
CLKBUF_X2 inst_17907 ( .A(net_17754), .Z(net_17755) );
CLKBUF_X2 inst_17094 ( .A(net_16941), .Z(net_16942) );
SDFF_X2 inst_1779 ( .D(net_7269), .SI(net_6966), .Q(net_6966), .SE(net_6283), .CK(net_14132) );
CLKBUF_X2 inst_19025 ( .A(net_18872), .Z(net_18873) );
DFFR_X2 inst_7299 ( .D(net_293), .QN(net_152), .CK(net_11607), .RN(x6501) );
SDFFR_X2 inst_2115 ( .SI(net_7173), .Q(net_7173), .D(net_4401), .SE(net_4362), .CK(net_17952), .RN(x6501) );
CLKBUF_X2 inst_18638 ( .A(net_18485), .Z(net_18486) );
CLKBUF_X2 inst_15910 ( .A(net_15757), .Z(net_15758) );
SDFF_X2 inst_1728 ( .Q(net_8187), .D(net_8187), .SI(net_2658), .SE(net_2561), .CK(net_15486) );
XNOR2_X2 inst_112 ( .B(net_7162), .ZN(net_4625), .A(net_4624) );
NOR3_X4 inst_3251 ( .A1(net_6128), .A2(net_2840), .ZN(net_2534), .A3(net_2453) );
CLKBUF_X2 inst_11161 ( .A(net_11008), .Z(net_11009) );
CLKBUF_X2 inst_9824 ( .A(net_9671), .Z(net_9672) );
CLKBUF_X2 inst_9523 ( .A(net_9370), .Z(net_9371) );
DFFR_X1 inst_7441 ( .QN(net_8920), .D(net_4763), .CK(net_17322), .RN(x6501) );
AOI22_X2 inst_8376 ( .A1(net_8597), .B1(net_8412), .A2(net_3864), .B2(net_3863), .ZN(net_3672) );
SDFFR_X1 inst_2724 ( .SI(net_9035), .Q(net_9035), .D(net_7464), .SE(net_3208), .CK(net_10665), .RN(x6501) );
CLKBUF_X2 inst_9353 ( .A(x12768), .Z(net_9201) );
DFFR_X2 inst_7067 ( .QN(net_7414), .D(net_4209), .CK(net_12308), .RN(x6501) );
CLKBUF_X2 inst_11334 ( .A(net_11181), .Z(net_11182) );
CLKBUF_X2 inst_12010 ( .A(net_11857), .Z(net_11858) );
INV_X4 inst_5751 ( .A(net_8944), .ZN(net_841) );
AOI22_X2 inst_8062 ( .B1(net_8173), .A1(net_7731), .B2(net_6101), .A2(net_6095), .ZN(net_4080) );
CLKBUF_X2 inst_10213 ( .A(net_9347), .Z(net_10061) );
SDFF_X2 inst_382 ( .SI(net_8395), .Q(net_8395), .SE(net_3969), .D(net_3955), .CK(net_13297) );
CLKBUF_X2 inst_9387 ( .A(net_9234), .Z(net_9235) );
SDFFR_X2 inst_2329 ( .SE(net_2260), .Q(net_330), .D(net_330), .CK(net_11506), .RN(x6501), .SI(x2633) );
CLKBUF_X2 inst_18294 ( .A(net_15385), .Z(net_18142) );
INV_X4 inst_6101 ( .ZN(net_486), .A(net_385) );
DFFR_X2 inst_7161 ( .QN(net_7206), .D(net_2771), .CK(net_15201), .RN(x6501) );
CLKBUF_X2 inst_10361 ( .A(net_9621), .Z(net_10209) );
CLKBUF_X2 inst_17548 ( .A(net_17395), .Z(net_17396) );
INV_X4 inst_6067 ( .A(net_8908), .ZN(net_5029) );
CLKBUF_X2 inst_10560 ( .A(net_10407), .Z(net_10408) );
CLKBUF_X2 inst_15040 ( .A(net_14887), .Z(net_14888) );
SDFF_X2 inst_1049 ( .SI(net_7310), .Q(net_6684), .D(net_6684), .SE(net_3126), .CK(net_11893) );
AOI22_X2 inst_8418 ( .B1(net_6652), .A1(net_6619), .A2(net_6213), .B2(net_6138), .ZN(net_3524) );
INV_X4 inst_5116 ( .A(net_8222), .ZN(net_4853) );
CLKBUF_X2 inst_17421 ( .A(net_17268), .Z(net_17269) );
AOI22_X2 inst_8085 ( .B1(net_8142), .A1(net_7904), .A2(net_6098), .ZN(net_6050), .B2(net_4190) );
NAND2_X2 inst_4575 ( .A2(net_2996), .ZN(net_2994), .A1(net_2993) );
CLKBUF_X2 inst_17085 ( .A(net_16301), .Z(net_16933) );
INV_X4 inst_6037 ( .A(net_8968), .ZN(net_1536) );
CLKBUF_X2 inst_13819 ( .A(net_11188), .Z(net_13667) );
CLKBUF_X2 inst_10547 ( .A(net_10394), .Z(net_10395) );
INV_X4 inst_5613 ( .A(net_6404), .ZN(net_1513) );
CLKBUF_X2 inst_12258 ( .A(net_11517), .Z(net_12106) );
CLKBUF_X2 inst_18749 ( .A(net_18596), .Z(net_18597) );
CLKBUF_X2 inst_9643 ( .A(net_9490), .Z(net_9491) );
CLKBUF_X2 inst_15113 ( .A(net_12769), .Z(net_14961) );
SDFF_X2 inst_580 ( .Q(net_8846), .D(net_8846), .SE(net_3964), .SI(net_3951), .CK(net_13418) );
CLKBUF_X2 inst_9249 ( .A(net_9096), .Z(net_9097) );
CLKBUF_X2 inst_13533 ( .A(net_13380), .Z(net_13381) );
CLKBUF_X2 inst_16519 ( .A(net_16366), .Z(net_16367) );
CLKBUF_X2 inst_16384 ( .A(net_16231), .Z(net_16232) );
CLKBUF_X2 inst_18217 ( .A(net_17266), .Z(net_18065) );
DFFR_X2 inst_7336 ( .Q(net_7342), .CK(net_11722), .D(x12891), .RN(x6501) );
CLKBUF_X2 inst_12647 ( .A(net_12494), .Z(net_12495) );
CLKBUF_X2 inst_11304 ( .A(net_11151), .Z(net_11152) );
CLKBUF_X2 inst_18128 ( .A(net_17975), .Z(net_17976) );
NOR2_X2 inst_3616 ( .A2(net_7427), .A1(net_7426), .ZN(net_2661) );
AOI221_X2 inst_8746 ( .B2(net_5657), .ZN(net_5653), .C2(net_5609), .A(net_5531), .B1(net_2724), .C1(net_363) );
AND2_X4 inst_9103 ( .ZN(net_2241), .A1(net_2123), .A2(net_2122) );
CLKBUF_X2 inst_13842 ( .A(net_13471), .Z(net_13690) );
SDFFR_X1 inst_2692 ( .SI(net_7553), .SE(net_5043), .CK(net_12739), .RN(x6501), .Q(x3874), .D(x3874) );
CLKBUF_X2 inst_17101 ( .A(net_16948), .Z(net_16949) );
CLKBUF_X2 inst_13580 ( .A(net_13427), .Z(net_13428) );
SDFF_X2 inst_1599 ( .Q(net_8134), .D(net_8134), .SI(net_2712), .SE(net_2541), .CK(net_17138) );
NOR2_X2 inst_3565 ( .ZN(net_1278), .A2(net_1152), .A1(net_760) );
INV_X8 inst_5026 ( .ZN(net_3984), .A(net_3319) );
DFFR_X2 inst_7348 ( .Q(net_7316), .CK(net_11382), .D(x13134), .RN(x6501) );
AOI22_X2 inst_8055 ( .B1(net_8172), .A1(net_7730), .B2(net_6101), .A2(net_6095), .ZN(net_4086) );
CLKBUF_X2 inst_14141 ( .A(net_13988), .Z(net_13989) );
INV_X4 inst_5687 ( .ZN(net_573), .A(net_148) );
AOI22_X2 inst_7922 ( .A1(net_8990), .A2(net_5456), .B2(net_5260), .ZN(net_4460), .B1(net_4459) );
CLKBUF_X2 inst_18744 ( .A(net_18591), .Z(net_18592) );
DFFS_X1 inst_6960 ( .D(net_2586), .CK(net_16569), .SN(x6501), .Q(x690) );
NAND3_X2 inst_3977 ( .ZN(net_2087), .A3(net_1796), .A2(net_1242), .A1(net_934) );
AOI222_X1 inst_8629 ( .B2(net_8238), .B1(net_4891), .C2(net_4889), .A1(net_4803), .ZN(net_4789), .C1(net_4457), .A2(net_3223) );
SDFFR_X2 inst_2593 ( .D(net_7380), .QN(net_7240), .SI(net_1943), .SE(net_1379), .CK(net_17515), .RN(x6501) );
CLKBUF_X2 inst_11717 ( .A(net_9513), .Z(net_11565) );
INV_X8 inst_5021 ( .ZN(net_5260), .A(net_4559) );
CLKBUF_X2 inst_9850 ( .A(net_9118), .Z(net_9698) );
CLKBUF_X2 inst_13550 ( .A(net_9686), .Z(net_13398) );
XNOR2_X2 inst_318 ( .ZN(net_946), .A(net_945), .B(net_193) );
CLKBUF_X2 inst_18055 ( .A(net_17902), .Z(net_17903) );
NAND2_X2 inst_4065 ( .ZN(net_5874), .A2(net_5770), .A1(net_3988) );
SDFF_X2 inst_1486 ( .SI(net_7291), .Q(net_7068), .D(net_7068), .SE(net_6280), .CK(net_15347) );
CLKBUF_X2 inst_13790 ( .A(net_10943), .Z(net_13638) );
SDFFR_X2 inst_2281 ( .SI(net_7394), .SE(net_2789), .Q(net_253), .D(net_253), .CK(net_17756), .RN(x6501) );
CLKBUF_X2 inst_13449 ( .A(net_13296), .Z(net_13297) );
SDFF_X2 inst_1175 ( .D(net_7340), .SI(net_6549), .Q(net_6549), .SE(net_3086), .CK(net_11856) );
CLKBUF_X2 inst_12666 ( .A(net_12513), .Z(net_12514) );
CLKBUF_X2 inst_13929 ( .A(net_11175), .Z(net_13777) );
CLKBUF_X2 inst_16778 ( .A(net_10749), .Z(net_16626) );
INV_X4 inst_5877 ( .A(net_8918), .ZN(net_2594) );
INV_X4 inst_5256 ( .ZN(net_2063), .A(net_1871) );
CLKBUF_X2 inst_12164 ( .A(net_12011), .Z(net_12012) );
CLKBUF_X2 inst_12208 ( .A(net_10251), .Z(net_12056) );
AOI22_X2 inst_8305 ( .B1(net_8733), .A1(net_8511), .B2(net_4350), .A2(net_4349), .ZN(net_3740) );
NAND2_X2 inst_4509 ( .A2(net_6209), .ZN(net_4321), .A1(net_1588) );
AOI21_X2 inst_8962 ( .ZN(net_3543), .B1(net_3542), .B2(net_3312), .A(net_2863) );
SDFF_X2 inst_395 ( .SI(net_8297), .Q(net_8297), .SE(net_3978), .D(net_3961), .CK(net_13214) );
CLKBUF_X2 inst_17634 ( .A(net_17481), .Z(net_17482) );
SDFF_X2 inst_841 ( .SI(net_8652), .Q(net_8652), .D(net_3963), .SE(net_3885), .CK(net_10058) );
CLKBUF_X2 inst_14106 ( .A(net_13953), .Z(net_13954) );
NAND3_X2 inst_3963 ( .ZN(net_2664), .A1(net_2384), .A2(net_1907), .A3(net_1906) );
DFFR_X2 inst_7328 ( .D(net_8286), .QN(net_8282), .CK(net_9971), .RN(x6501) );
CLKBUF_X2 inst_13682 ( .A(net_13529), .Z(net_13530) );
CLKBUF_X2 inst_13412 ( .A(net_13259), .Z(net_13260) );
NAND2_X2 inst_4895 ( .A2(net_7377), .ZN(net_650), .A1(net_166) );
INV_X2 inst_6361 ( .ZN(net_2166), .A(net_2072) );
CLKBUF_X2 inst_13538 ( .A(net_13385), .Z(net_13386) );
CLKBUF_X2 inst_17457 ( .A(net_17304), .Z(net_17305) );
NAND3_X2 inst_3896 ( .ZN(net_5642), .A1(net_5571), .A3(net_5505), .A2(net_5410) );
NAND4_X2 inst_3679 ( .A4(net_6030), .A1(net_6029), .ZN(net_4586), .A2(net_4016), .A3(net_4015) );
SDFF_X2 inst_1558 ( .Q(net_7882), .D(net_7882), .SI(net_2702), .SE(net_2543), .CK(net_18053) );
CLKBUF_X2 inst_14212 ( .A(net_14059), .Z(net_14060) );
OAI33_X1 inst_2906 ( .B3(net_9010), .B2(net_6169), .ZN(net_2430), .B1(net_2429), .A3(net_2429), .A1(net_2186), .A2(net_722) );
INV_X4 inst_5848 ( .A(net_7509), .ZN(net_3239) );
CLKBUF_X2 inst_14622 ( .A(net_14469), .Z(net_14470) );
CLKBUF_X2 inst_13398 ( .A(net_13245), .Z(net_13246) );
CLKBUF_X2 inst_14206 ( .A(net_14053), .Z(net_14054) );
NAND3_X2 inst_3886 ( .ZN(net_5853), .A3(net_5852), .A1(net_5751), .A2(net_1315) );
CLKBUF_X2 inst_12836 ( .A(net_12683), .Z(net_12684) );
AOI221_X2 inst_8797 ( .C2(net_6187), .B2(net_5609), .A(net_4898), .ZN(net_4880), .B1(net_368), .C1(net_192) );
AND2_X4 inst_9072 ( .ZN(net_6104), .A2(net_3248), .A1(net_3215) );
CLKBUF_X2 inst_13201 ( .A(net_10700), .Z(net_13049) );
CLKBUF_X2 inst_9505 ( .A(net_9090), .Z(net_9353) );
CLKBUF_X2 inst_11692 ( .A(net_10356), .Z(net_11540) );
CLKBUF_X2 inst_10643 ( .A(net_10490), .Z(net_10491) );
CLKBUF_X2 inst_11510 ( .A(net_9768), .Z(net_11358) );
CLKBUF_X2 inst_9890 ( .A(net_9737), .Z(net_9738) );
CLKBUF_X2 inst_12127 ( .A(net_11974), .Z(net_11975) );
SDFF_X2 inst_920 ( .SI(net_8707), .Q(net_8707), .SE(net_6195), .D(net_3977), .CK(net_13023) );
NOR2_X2 inst_3454 ( .A1(net_3023), .ZN(net_2918), .A2(net_2813) );
INV_X2 inst_6298 ( .ZN(net_4200), .A(net_3909) );
CLKBUF_X2 inst_18010 ( .A(net_17857), .Z(net_17858) );
INV_X4 inst_5741 ( .A(net_8281), .ZN(net_958) );
INV_X2 inst_6571 ( .ZN(net_888), .A(net_207) );
CLKBUF_X2 inst_16903 ( .A(net_16750), .Z(net_16751) );
INV_X4 inst_6116 ( .A(net_7481), .ZN(net_1658) );
CLKBUF_X2 inst_11629 ( .A(net_9655), .Z(net_11477) );
CLKBUF_X2 inst_13797 ( .A(net_13644), .Z(net_13645) );
OR2_X2 inst_2889 ( .ZN(net_1710), .A1(net_1685), .A2(net_1577) );
CLKBUF_X2 inst_14203 ( .A(net_14050), .Z(net_14051) );
CLKBUF_X2 inst_18839 ( .A(net_18686), .Z(net_18687) );
CLKBUF_X2 inst_16935 ( .A(net_16782), .Z(net_16783) );
CLKBUF_X2 inst_10109 ( .A(net_9956), .Z(net_9957) );
CLKBUF_X2 inst_11380 ( .A(net_11227), .Z(net_11228) );
CLKBUF_X2 inst_15265 ( .A(net_15112), .Z(net_15113) );
AOI22_X2 inst_8034 ( .B1(net_8033), .A1(net_7999), .B2(net_6102), .A2(net_6097), .ZN(net_4104) );
CLKBUF_X2 inst_13743 ( .A(net_13590), .Z(net_13591) );
SDFFR_X2 inst_2189 ( .SI(net_8965), .Q(net_8965), .SE(net_2967), .D(net_2012), .CK(net_17580), .RN(x6501) );
INV_X4 inst_5448 ( .A(net_881), .ZN(net_811) );
XNOR2_X2 inst_315 ( .A(net_7586), .B(net_3390), .ZN(net_950) );
NAND2_X2 inst_4198 ( .ZN(net_5300), .A2(net_5178), .A1(net_5057) );
CLKBUF_X2 inst_13176 ( .A(net_11187), .Z(net_13024) );
CLKBUF_X2 inst_14989 ( .A(net_14836), .Z(net_14837) );
XNOR2_X2 inst_216 ( .B(net_8894), .ZN(net_1424), .A(net_1423) );
AOI21_X2 inst_8992 ( .ZN(net_1495), .B1(net_1494), .A(net_1353), .B2(net_1141) );
CLKBUF_X2 inst_16708 ( .A(net_16555), .Z(net_16556) );
CLKBUF_X2 inst_15126 ( .A(net_14973), .Z(net_14974) );
CLKBUF_X2 inst_14858 ( .A(net_10087), .Z(net_14706) );
CLKBUF_X2 inst_13099 ( .A(net_12946), .Z(net_12947) );
SDFFS_X2 inst_2060 ( .SI(net_8289), .Q(net_8289), .SE(net_3552), .D(net_959), .CK(net_11194), .SN(x6501) );
CLKBUF_X2 inst_12987 ( .A(net_10355), .Z(net_12835) );
SDFFR_X1 inst_2680 ( .SI(net_7538), .SE(net_5043), .CK(net_9699), .RN(x6501), .Q(x4082), .D(x4082) );
AOI221_X2 inst_8771 ( .C1(net_8987), .B2(net_5538), .C2(net_5456), .ZN(net_5277), .A(net_4873), .B1(net_416) );
DFFR_X2 inst_7321 ( .D(net_8287), .QN(net_8283), .CK(net_9975), .RN(x6501) );
CLKBUF_X2 inst_9225 ( .A(net_9072), .Z(net_9073) );
SDFF_X2 inst_1795 ( .D(net_7282), .SI(net_6979), .Q(net_6979), .SE(net_6283), .CK(net_16201) );
SDFF_X2 inst_828 ( .SI(net_8488), .Q(net_8488), .D(net_3947), .SE(net_3884), .CK(net_12419) );
NAND2_X2 inst_4697 ( .A1(net_6411), .A2(net_1902), .ZN(net_1893) );
CLKBUF_X2 inst_18173 ( .A(net_14147), .Z(net_18021) );
CLKBUF_X2 inst_13522 ( .A(net_13369), .Z(net_13370) );
DFFR_X2 inst_7218 ( .D(net_2359), .QN(net_221), .CK(net_17467), .RN(x6501) );
CLKBUF_X2 inst_17072 ( .A(net_16919), .Z(net_16920) );
NAND2_X2 inst_4164 ( .ZN(net_5348), .A1(net_5092), .A2(net_5091) );
CLKBUF_X2 inst_15852 ( .A(net_15699), .Z(net_15700) );
CLKBUF_X2 inst_16446 ( .A(net_11106), .Z(net_16294) );
CLKBUF_X2 inst_17540 ( .A(net_17387), .Z(net_17388) );
AOI21_X2 inst_8899 ( .B2(net_5871), .ZN(net_5781), .A(net_5758), .B1(x186) );
CLKBUF_X2 inst_13919 ( .A(net_13766), .Z(net_13767) );
AOI22_X2 inst_8052 ( .B1(net_8036), .A1(net_8002), .B2(net_6102), .A2(net_6097), .ZN(net_4089) );
CLKBUF_X2 inst_10854 ( .A(net_10701), .Z(net_10702) );
CLKBUF_X2 inst_17766 ( .A(net_17613), .Z(net_17614) );
INV_X2 inst_6182 ( .ZN(net_5847), .A(net_5792) );
DFFR_X1 inst_7382 ( .D(net_5919), .CK(net_17186), .RN(x6501), .Q(x208) );
AOI221_X2 inst_8749 ( .B2(net_5657), .C2(net_5609), .ZN(net_5608), .A(net_5516), .B1(net_2735), .C1(net_365) );
INV_X2 inst_6240 ( .ZN(net_4896), .A(net_4801) );
CLKBUF_X2 inst_9629 ( .A(net_9476), .Z(net_9477) );
CLKBUF_X2 inst_11426 ( .A(net_11273), .Z(net_11274) );
CLKBUF_X2 inst_10127 ( .A(net_9974), .Z(net_9975) );
AND2_X4 inst_9137 ( .ZN(net_1383), .A2(net_798), .A1(net_174) );
CLKBUF_X2 inst_10794 ( .A(net_10233), .Z(net_10642) );
CLKBUF_X2 inst_10951 ( .A(net_10798), .Z(net_10799) );
OAI21_X2 inst_3050 ( .B2(net_8231), .B1(net_4850), .ZN(net_4761), .A(net_2627) );
CLKBUF_X2 inst_11349 ( .A(net_11041), .Z(net_11197) );
CLKBUF_X2 inst_13916 ( .A(net_13763), .Z(net_13764) );
AOI22_X2 inst_8491 ( .B1(net_6612), .A1(net_6579), .A2(net_6257), .B2(net_6110), .ZN(net_3449) );
CLKBUF_X2 inst_18276 ( .A(net_18123), .Z(net_18124) );
NAND3_X2 inst_3913 ( .ZN(net_5625), .A1(net_5554), .A3(net_5488), .A2(net_5342) );
CLKBUF_X2 inst_19137 ( .A(net_10634), .Z(net_18985) );
INV_X4 inst_5807 ( .A(net_6285), .ZN(net_2512) );
CLKBUF_X2 inst_12625 ( .A(net_12472), .Z(net_12473) );
DFFR_X1 inst_7484 ( .QN(net_7430), .D(net_4205), .CK(net_12380), .RN(x6501) );
SDFF_X2 inst_1941 ( .SI(net_8074), .Q(net_8074), .D(net_2704), .SE(net_2508), .CK(net_16970) );
INV_X2 inst_6247 ( .ZN(net_4859), .A(net_4753) );
XOR2_X2 inst_9 ( .A(net_2993), .Z(net_2029), .B(net_1696) );
NOR2_X2 inst_3358 ( .ZN(net_5567), .A1(net_5396), .A2(net_5395) );
DFF_X1 inst_6719 ( .Q(net_6765), .D(net_5650), .CK(net_9275) );
CLKBUF_X2 inst_18751 ( .A(net_18598), .Z(net_18599) );
SDFF_X2 inst_1594 ( .Q(net_8126), .D(net_8126), .SI(net_2589), .SE(net_2541), .CK(net_18861) );
SDFF_X2 inst_902 ( .SI(net_8719), .Q(net_8719), .SE(net_6195), .D(net_3973), .CK(net_13158) );
CLKBUF_X2 inst_15810 ( .A(net_12539), .Z(net_15658) );
NOR2_X2 inst_3489 ( .ZN(net_2092), .A1(net_2091), .A2(net_1741) );
CLKBUF_X2 inst_12224 ( .A(net_12071), .Z(net_12072) );
SDFF_X2 inst_778 ( .SI(net_8346), .Q(net_8346), .D(net_3945), .SE(net_3880), .CK(net_13096) );
CLKBUF_X2 inst_10118 ( .A(net_9718), .Z(net_9966) );
CLKBUF_X2 inst_16581 ( .A(net_14091), .Z(net_16429) );
CLKBUF_X2 inst_17405 ( .A(net_11384), .Z(net_17253) );
AOI22_X2 inst_7912 ( .B1(net_7516), .B2(net_5260), .ZN(net_4502), .A2(net_4501), .A1(net_2739) );
CLKBUF_X2 inst_14842 ( .A(net_14689), .Z(net_14690) );
CLKBUF_X2 inst_11486 ( .A(net_10178), .Z(net_11334) );
AOI22_X2 inst_7810 ( .A2(net_8219), .B2(net_6144), .A1(net_4764), .ZN(net_4754), .B1(net_4732) );
AOI221_X2 inst_8845 ( .B1(net_8556), .C1(net_8445), .C2(net_6263), .B2(net_6262), .ZN(net_6239), .A(net_4267) );
CLKBUF_X2 inst_17945 ( .A(net_16679), .Z(net_17793) );
AOI22_X2 inst_8353 ( .A1(net_8627), .B1(net_8442), .A2(net_3864), .B2(net_3863), .ZN(net_3695) );
CLKBUF_X2 inst_12855 ( .A(net_12702), .Z(net_12703) );
CLKBUF_X2 inst_13895 ( .A(net_11483), .Z(net_13743) );
SDFF_X2 inst_781 ( .SI(net_8350), .Q(net_8350), .D(net_3944), .SE(net_3880), .CK(net_10824) );
CLKBUF_X2 inst_18034 ( .A(net_17881), .Z(net_17882) );
CLKBUF_X2 inst_12033 ( .A(net_11880), .Z(net_11881) );
NAND2_X4 inst_4042 ( .ZN(net_6258), .A1(net_6251), .A2(net_2210) );
CLKBUF_X2 inst_12368 ( .A(net_12215), .Z(net_12216) );
CLKBUF_X2 inst_13409 ( .A(net_9073), .Z(net_13257) );
NAND4_X2 inst_3696 ( .A4(net_6224), .A1(net_6223), .ZN(net_4441), .A2(net_3786), .A3(net_3785) );
CLKBUF_X2 inst_9450 ( .A(net_9059), .Z(net_9298) );
CLKBUF_X2 inst_17593 ( .A(net_17440), .Z(net_17441) );
CLKBUF_X2 inst_18731 ( .A(net_18578), .Z(net_18579) );
CLKBUF_X2 inst_9971 ( .A(net_9818), .Z(net_9819) );
CLKBUF_X2 inst_16883 ( .A(net_16730), .Z(net_16731) );
DFFR_X2 inst_7053 ( .Q(net_7511), .D(net_4831), .CK(net_17638), .RN(x6501) );
SDFF_X2 inst_1928 ( .SI(net_8055), .Q(net_8055), .D(net_2706), .SE(net_2508), .CK(net_15230) );
SDFF_X2 inst_1967 ( .D(net_7276), .SI(net_7013), .Q(net_7013), .SE(net_6277), .CK(net_17335) );
NAND2_X2 inst_4485 ( .A2(net_5267), .ZN(net_4493), .A1(net_170) );
CLKBUF_X2 inst_13733 ( .A(net_13580), .Z(net_13581) );
CLKBUF_X2 inst_12944 ( .A(net_12791), .Z(net_12792) );
SDFF_X2 inst_1947 ( .SI(net_8051), .Q(net_8051), .D(net_2658), .SE(net_2508), .CK(net_15228) );
CLKBUF_X2 inst_10967 ( .A(net_9692), .Z(net_10815) );
DFFR_X2 inst_7318 ( .D(net_6826), .QN(net_6823), .CK(net_15089), .RN(x6501) );
AOI22_X2 inst_8030 ( .B1(net_8101), .A1(net_7761), .B2(net_6108), .A2(net_6096), .ZN(net_4108) );
INV_X2 inst_6285 ( .ZN(net_4215), .A(net_3924) );
CLKBUF_X2 inst_18186 ( .A(net_18033), .Z(net_18034) );
NAND2_X2 inst_4585 ( .ZN(net_3149), .A2(net_2908), .A1(net_2216) );
AOI22_X2 inst_8105 ( .B1(net_8077), .A1(net_7873), .B2(net_6107), .ZN(net_5994), .A2(net_4400) );
CLKBUF_X2 inst_15143 ( .A(net_14990), .Z(net_14991) );
CLKBUF_X2 inst_18102 ( .A(net_17949), .Z(net_17950) );
AND2_X4 inst_9126 ( .ZN(net_1425), .A2(net_905), .A1(net_185) );
CLKBUF_X2 inst_9539 ( .A(net_9386), .Z(net_9387) );
CLKBUF_X2 inst_19141 ( .A(net_18667), .Z(net_18989) );
CLKBUF_X2 inst_15304 ( .A(net_15151), .Z(net_15152) );
CLKBUF_X2 inst_11294 ( .A(net_10561), .Z(net_11142) );
DFFR_X1 inst_7573 ( .Q(net_7627), .D(net_7624), .CK(net_18011), .RN(x6501) );
CLKBUF_X2 inst_16830 ( .A(net_16677), .Z(net_16678) );
SDFF_X2 inst_659 ( .Q(net_8432), .D(net_8432), .SI(net_3955), .SE(net_3934), .CK(net_13254) );
CLKBUF_X2 inst_17194 ( .A(net_17041), .Z(net_17042) );
DFFS_X2 inst_6890 ( .QN(net_6753), .D(net_2895), .CK(net_9120), .SN(x6501) );
CLKBUF_X2 inst_11747 ( .A(net_11594), .Z(net_11595) );
CLKBUF_X2 inst_12868 ( .A(net_9176), .Z(net_12716) );
CLKBUF_X2 inst_12883 ( .A(net_12730), .Z(net_12731) );
INV_X4 inst_5273 ( .ZN(net_2049), .A(net_1688) );
AOI22_X2 inst_8094 ( .B1(net_8041), .A1(net_8007), .B2(net_6102), .A2(net_6097), .ZN(net_4053) );
INV_X4 inst_5505 ( .A(net_3600), .ZN(net_693) );
CLKBUF_X2 inst_10289 ( .A(net_10136), .Z(net_10137) );
OAI211_X2 inst_3199 ( .ZN(net_3080), .C1(net_2530), .C2(net_2525), .B(net_2445), .A(net_2249) );
INV_X2 inst_6178 ( .ZN(net_5908), .A(net_5862) );
NOR2_X2 inst_3612 ( .A2(net_7518), .A1(net_7517), .ZN(net_1337) );
SDFF_X2 inst_1581 ( .Q(net_8033), .D(net_8033), .SI(net_2749), .SE(net_2545), .CK(net_16494) );
CLKBUF_X2 inst_17952 ( .A(net_17799), .Z(net_17800) );
SDFFR_X2 inst_2312 ( .SE(net_2678), .D(net_1484), .SI(net_403), .Q(net_403), .CK(net_16665), .RN(x6501) );
INV_X4 inst_5336 ( .A(net_7212), .ZN(net_1507) );
NOR2_X2 inst_3500 ( .ZN(net_4513), .A2(net_1880), .A1(net_1311) );
CLKBUF_X2 inst_17248 ( .A(net_17095), .Z(net_17096) );
INV_X2 inst_6381 ( .A(net_1479), .ZN(net_1341) );
CLKBUF_X2 inst_10526 ( .A(net_9542), .Z(net_10374) );
DFFR_X2 inst_7103 ( .QN(net_9004), .D(net_3257), .CK(net_13459), .RN(x6501) );
SDFFR_X2 inst_2241 ( .Q(net_7455), .D(net_7455), .SE(net_2863), .CK(net_12915), .SI(x13541), .RN(x6501) );
CLKBUF_X2 inst_13419 ( .A(net_13266), .Z(net_13267) );
AOI22_X2 inst_8165 ( .B1(net_8815), .A1(net_8334), .A2(net_6265), .B2(net_6253), .ZN(net_6072) );
SDFFR_X2 inst_2182 ( .QN(net_7571), .D(net_3960), .SE(net_3144), .SI(net_595), .CK(net_10866), .RN(x6501) );
AOI22_X2 inst_8334 ( .B1(net_8588), .A1(net_8477), .A2(net_6263), .B2(net_6262), .ZN(net_3713) );
SDFFR_X1 inst_2667 ( .D(net_6764), .SE(net_4506), .CK(net_11531), .RN(x6501), .SI(x1935), .Q(x1935) );
CLKBUF_X2 inst_17049 ( .A(net_16896), .Z(net_16897) );
SDFF_X2 inst_987 ( .D(net_7324), .SI(net_6632), .Q(net_6632), .SE(net_3123), .CK(net_9873) );
NAND2_X2 inst_4194 ( .ZN(net_5305), .A1(net_5062), .A2(net_5061) );
CLKBUF_X2 inst_9376 ( .A(net_9223), .Z(net_9224) );
OAI21_X2 inst_3006 ( .ZN(net_5757), .A(net_5756), .B2(net_5755), .B1(net_518) );
CLKBUF_X2 inst_17026 ( .A(net_16873), .Z(net_16874) );
CLKBUF_X2 inst_9703 ( .A(net_9550), .Z(net_9551) );
CLKBUF_X2 inst_18044 ( .A(net_16002), .Z(net_17892) );
CLKBUF_X2 inst_15350 ( .A(net_10064), .Z(net_15198) );
SDFF_X2 inst_371 ( .SI(net_8298), .Q(net_8298), .SE(net_3978), .D(net_3943), .CK(net_13376) );
MUX2_X2 inst_4962 ( .A(net_7384), .S(net_2370), .Z(net_2361), .B(net_799) );
INV_X2 inst_6498 ( .A(net_9050), .ZN(net_903) );
CLKBUF_X2 inst_10768 ( .A(net_9130), .Z(net_10616) );
NAND2_X2 inst_4619 ( .A2(net_6144), .ZN(net_2603), .A1(net_2602) );
CLKBUF_X2 inst_18511 ( .A(net_18358), .Z(net_18359) );
CLKBUF_X2 inst_17301 ( .A(net_15991), .Z(net_17149) );
NAND4_X2 inst_3684 ( .ZN(net_4453), .A4(net_4352), .A1(net_3869), .A2(net_3868), .A3(net_3865) );
SDFF_X2 inst_628 ( .SI(net_8540), .Q(net_8540), .SE(net_3979), .D(net_3956), .CK(net_10925) );
DFFR_X1 inst_7470 ( .Q(net_7442), .D(net_4230), .CK(net_12935), .RN(x6501) );
NAND4_X2 inst_3642 ( .ZN(net_4942), .A1(net_4715), .A4(net_4561), .A3(net_4532), .A2(net_4479) );
CLKBUF_X2 inst_11873 ( .A(net_11720), .Z(net_11721) );
CLKBUF_X2 inst_17883 ( .A(net_17730), .Z(net_17731) );
OAI21_X2 inst_3092 ( .ZN(net_2862), .B2(net_2861), .A(net_1873), .B1(net_1709) );
INV_X2 inst_6587 ( .A(net_6113), .ZN(net_6112) );
CLKBUF_X2 inst_14162 ( .A(net_9118), .Z(net_14010) );
CLKBUF_X2 inst_17911 ( .A(net_17758), .Z(net_17759) );
NOR2_X2 inst_3395 ( .ZN(net_4564), .A2(net_4512), .A1(net_4394) );
SDFF_X2 inst_1130 ( .D(net_7337), .SI(net_6579), .Q(net_6579), .SE(net_3070), .CK(net_9453) );
CLKBUF_X2 inst_9300 ( .A(net_9091), .Z(net_9148) );
CLKBUF_X2 inst_18239 ( .A(net_10412), .Z(net_18087) );
CLKBUF_X2 inst_18617 ( .A(net_18464), .Z(net_18465) );
CLKBUF_X2 inst_18405 ( .A(net_18252), .Z(net_18253) );
INV_X2 inst_6304 ( .ZN(net_3900), .A(net_3602) );
CLKBUF_X2 inst_12706 ( .A(net_12553), .Z(net_12554) );
CLKBUF_X2 inst_17341 ( .A(net_17188), .Z(net_17189) );
AOI22_X2 inst_7851 ( .A2(net_5595), .ZN(net_4656), .B2(net_4388), .B1(net_2612), .A1(net_321) );
AOI21_X2 inst_8996 ( .B1(net_6414), .B2(net_6413), .ZN(net_1576), .A(net_1316) );
CLKBUF_X2 inst_15748 ( .A(net_15595), .Z(net_15596) );
CLKBUF_X2 inst_11823 ( .A(net_11670), .Z(net_11671) );
CLKBUF_X2 inst_18506 ( .A(net_18353), .Z(net_18354) );
INV_X4 inst_5425 ( .A(net_7305), .ZN(net_1494) );
CLKBUF_X2 inst_9304 ( .A(net_9071), .Z(net_9152) );
SDFF_X2 inst_1363 ( .SI(net_7263), .Q(net_7120), .D(net_7120), .SE(net_6279), .CK(net_17092) );
NAND2_X2 inst_4851 ( .A1(net_1243), .A2(net_955), .ZN(net_899) );
CLKBUF_X2 inst_18097 ( .A(net_17944), .Z(net_17945) );
CLKBUF_X2 inst_17038 ( .A(net_16885), .Z(net_16886) );
CLKBUF_X2 inst_17357 ( .A(net_14354), .Z(net_17205) );
AOI22_X2 inst_8059 ( .B1(net_8037), .A1(net_8003), .B2(net_6102), .A2(net_6097), .ZN(net_4083) );
CLKBUF_X2 inst_12388 ( .A(net_12235), .Z(net_12236) );
CLKBUF_X2 inst_11372 ( .A(net_11219), .Z(net_11220) );
CLKBUF_X2 inst_11806 ( .A(net_11653), .Z(net_11654) );
CLKBUF_X2 inst_11992 ( .A(net_11839), .Z(net_11840) );
CLKBUF_X2 inst_15736 ( .A(net_15583), .Z(net_15584) );
SDFFR_X2 inst_2127 ( .SI(net_7189), .Q(net_7189), .D(net_6440), .SE(net_4362), .CK(net_17838), .RN(x6501) );
HA_X1 inst_6688 ( .A(net_3111), .S(net_2977), .CO(net_2976), .B(net_2805) );
CLKBUF_X2 inst_13626 ( .A(net_13473), .Z(net_13474) );
CLKBUF_X2 inst_13689 ( .A(net_13536), .Z(net_13537) );
CLKBUF_X2 inst_10611 ( .A(net_10458), .Z(net_10459) );
CLKBUF_X2 inst_16974 ( .A(net_16821), .Z(net_16822) );
SDFFR_X2 inst_2268 ( .SI(net_7379), .SE(net_2793), .Q(net_238), .D(net_238), .CK(net_17833), .RN(x6501) );
SDFF_X2 inst_1373 ( .Q(net_8213), .D(net_8213), .SI(net_2703), .SE(net_2561), .CK(net_14022) );
SDFFR_X2 inst_2458 ( .QN(net_7478), .SE(net_3354), .SI(net_3128), .CK(net_12159), .D(x13353), .RN(x6501) );
DFFR_X2 inst_7285 ( .D(net_390), .Q(net_265), .CK(net_13522), .RN(x6501) );
AOI22_X2 inst_8474 ( .B1(net_6674), .A1(net_6641), .A2(net_6213), .B2(net_6138), .ZN(net_3466) );
CLKBUF_X2 inst_14303 ( .A(net_10290), .Z(net_14151) );
OAI21_X2 inst_3155 ( .B2(net_1984), .ZN(net_1978), .A(net_1977), .B1(net_1976) );
CLKBUF_X2 inst_9923 ( .A(net_9770), .Z(net_9771) );
OAI21_X2 inst_3134 ( .B2(net_2247), .A(net_2172), .ZN(net_2072), .B1(net_2071) );
INV_X4 inst_5481 ( .A(net_1150), .ZN(net_1075) );
NAND2_X4 inst_4043 ( .A1(net_2327), .ZN(net_2324), .A2(net_852) );
HA_X1 inst_6710 ( .CO(net_1570), .S(net_1238), .A(net_1237), .B(net_1236) );
CLKBUF_X2 inst_11787 ( .A(net_11634), .Z(net_11635) );
AOI22_X2 inst_8407 ( .B1(net_8564), .A1(net_8453), .A2(net_6263), .B2(net_6262), .ZN(net_3645) );
CLKBUF_X2 inst_18647 ( .A(net_18494), .Z(net_18495) );
CLKBUF_X2 inst_11999 ( .A(net_11846), .Z(net_11847) );
INV_X4 inst_5755 ( .ZN(net_561), .A(x2400) );
CLKBUF_X2 inst_11933 ( .A(net_11029), .Z(net_11781) );
CLKBUF_X2 inst_16163 ( .A(net_16010), .Z(net_16011) );
CLKBUF_X2 inst_17432 ( .A(net_17279), .Z(net_17280) );
AOI22_X2 inst_8122 ( .B1(net_8116), .A1(net_7878), .A2(net_6098), .B2(net_4190), .ZN(net_4027) );
CLKBUF_X2 inst_17620 ( .A(net_9340), .Z(net_17468) );
CLKBUF_X2 inst_15077 ( .A(net_14924), .Z(net_14925) );
CLKBUF_X2 inst_13435 ( .A(net_11597), .Z(net_13283) );
CLKBUF_X2 inst_15728 ( .A(net_12716), .Z(net_15576) );
CLKBUF_X2 inst_12349 ( .A(net_12196), .Z(net_12197) );
CLKBUF_X2 inst_12490 ( .A(net_9651), .Z(net_12338) );
NAND2_X2 inst_4588 ( .A1(net_7353), .ZN(net_2883), .A2(net_2881) );
CLKBUF_X2 inst_12755 ( .A(net_10804), .Z(net_12603) );
CLKBUF_X2 inst_13746 ( .A(net_11466), .Z(net_13594) );
AND2_X4 inst_9099 ( .ZN(net_5027), .A1(net_2262), .A2(net_2090) );
NAND2_X4 inst_4049 ( .ZN(net_2461), .A2(net_2299), .A1(net_1695) );
SDFFR_X1 inst_2702 ( .SI(net_7534), .SE(net_5043), .CK(net_11930), .RN(x6501), .Q(x4132), .D(x4132) );
INV_X4 inst_5067 ( .ZN(net_5883), .A(net_5845) );
CLKBUF_X2 inst_15063 ( .A(net_14910), .Z(net_14911) );
CLKBUF_X2 inst_12820 ( .A(net_10605), .Z(net_12668) );
OAI22_X2 inst_2910 ( .A2(net_8232), .B2(net_6133), .A1(net_4954), .ZN(net_4874), .B1(net_1417) );
NAND2_X2 inst_4670 ( .ZN(net_2396), .A2(net_2162), .A1(net_1473) );
INV_X4 inst_5701 ( .A(net_7518), .ZN(net_2569) );
CLKBUF_X2 inst_15178 ( .A(net_15025), .Z(net_15026) );
CLKBUF_X2 inst_16586 ( .A(net_14945), .Z(net_16434) );
XNOR2_X2 inst_145 ( .ZN(net_2228), .B(net_2141), .A(net_2140) );
CLKBUF_X2 inst_13703 ( .A(net_11733), .Z(net_13551) );
NAND2_X2 inst_4594 ( .ZN(net_3064), .A1(net_2835), .A2(net_2834) );
INV_X4 inst_5355 ( .A(net_2556), .ZN(net_1155) );
CLKBUF_X2 inst_9689 ( .A(net_9536), .Z(net_9537) );
CLKBUF_X2 inst_15223 ( .A(net_15070), .Z(net_15071) );
INV_X2 inst_6214 ( .ZN(net_5496), .A(net_5373) );
CLKBUF_X2 inst_10199 ( .A(net_10046), .Z(net_10047) );
CLKBUF_X2 inst_17338 ( .A(net_17185), .Z(net_17186) );
SDFF_X2 inst_1437 ( .SI(net_7280), .Q(net_7097), .D(net_7097), .SE(net_6278), .CK(net_19037) );
INV_X4 inst_5345 ( .ZN(net_2946), .A(net_2531) );
CLKBUF_X2 inst_12240 ( .A(net_9284), .Z(net_12088) );
CLKBUF_X2 inst_18006 ( .A(net_17853), .Z(net_17854) );
CLKBUF_X2 inst_17483 ( .A(net_17330), .Z(net_17331) );
AND2_X4 inst_9119 ( .A2(net_8217), .ZN(net_2261), .A1(net_1082) );
CLKBUF_X2 inst_9292 ( .A(net_9098), .Z(net_9140) );
CLKBUF_X2 inst_10557 ( .A(net_10404), .Z(net_10405) );
CLKBUF_X2 inst_13661 ( .A(net_13508), .Z(net_13509) );
SDFFR_X2 inst_2533 ( .QN(net_6373), .D(net_2148), .SE(net_2147), .SI(net_1954), .CK(net_18149), .RN(x6501) );
XOR2_X2 inst_27 ( .Z(net_1228), .A(net_596), .B(net_195) );
AOI221_X2 inst_8790 ( .B2(net_5595), .ZN(net_4911), .C2(net_4881), .A(net_4639), .B1(net_330), .C1(net_248) );
CLKBUF_X2 inst_10741 ( .A(net_10588), .Z(net_10589) );
NAND2_X2 inst_4446 ( .A1(net_6846), .A2(net_5016), .ZN(net_4981) );
CLKBUF_X2 inst_14849 ( .A(net_13145), .Z(net_14697) );
CLKBUF_X2 inst_16721 ( .A(net_16568), .Z(net_16569) );
CLKBUF_X2 inst_11761 ( .A(net_11608), .Z(net_11609) );
CLKBUF_X2 inst_10063 ( .A(net_9910), .Z(net_9911) );
CLKBUF_X2 inst_16060 ( .A(net_15907), .Z(net_15908) );
CLKBUF_X2 inst_15397 ( .A(net_15244), .Z(net_15245) );
CLKBUF_X2 inst_15807 ( .A(net_15654), .Z(net_15655) );
INV_X2 inst_6420 ( .A(net_948), .ZN(net_770) );
CLKBUF_X2 inst_15879 ( .A(net_15726), .Z(net_15727) );
INV_X4 inst_5230 ( .ZN(net_5746), .A(net_2252) );
SDFF_X2 inst_639 ( .SI(net_8554), .Q(net_8554), .SE(net_3979), .D(net_3949), .CK(net_12792) );
AND3_X4 inst_9045 ( .ZN(net_1654), .A3(net_154), .A2(net_153), .A1(net_152) );
CLKBUF_X2 inst_14687 ( .A(net_14534), .Z(net_14535) );
NAND3_X2 inst_3939 ( .ZN(net_4920), .A3(net_4679), .A1(net_4668), .A2(net_4644) );
CLKBUF_X2 inst_19095 ( .A(net_17446), .Z(net_18943) );
CLKBUF_X2 inst_17819 ( .A(net_17666), .Z(net_17667) );
SDFFR_X2 inst_2167 ( .QN(net_7591), .D(net_3940), .SE(net_3144), .SI(net_547), .CK(net_10392), .RN(x6501) );
DFFR_X2 inst_7008 ( .QN(net_6315), .D(net_5787), .CK(net_16943), .RN(x6501) );
CLKBUF_X2 inst_12193 ( .A(net_12040), .Z(net_12041) );
DFFR_X1 inst_7412 ( .D(net_5735), .Q(net_257), .CK(net_17489), .RN(x6501) );
INV_X2 inst_6328 ( .ZN(net_3213), .A(net_3183) );
SDFF_X2 inst_1651 ( .SI(net_7706), .Q(net_7706), .D(net_2705), .SE(net_2559), .CK(net_18543) );
NAND2_X2 inst_4248 ( .A1(net_7027), .A2(net_5249), .ZN(net_5212) );
CLKBUF_X2 inst_12561 ( .A(net_11469), .Z(net_12409) );
CLKBUF_X2 inst_12176 ( .A(net_12023), .Z(net_12024) );
AOI22_X2 inst_8281 ( .B1(net_8581), .A1(net_8470), .A2(net_6263), .B2(net_6262), .ZN(net_3760) );
CLKBUF_X2 inst_9758 ( .A(net_9180), .Z(net_9606) );
CLKBUF_X2 inst_15695 ( .A(net_15542), .Z(net_15543) );
INV_X2 inst_6451 ( .A(net_7430), .ZN(net_591) );
CLKBUF_X2 inst_11159 ( .A(net_10488), .Z(net_11007) );
SDFF_X2 inst_1137 ( .D(net_7315), .SI(net_6557), .Q(net_6557), .SE(net_3070), .CK(net_9913) );
CLKBUF_X2 inst_15254 ( .A(net_13604), .Z(net_15102) );
SDFF_X2 inst_1389 ( .SI(net_7731), .Q(net_7731), .D(net_2639), .SE(net_2559), .CK(net_17147) );
CLKBUF_X2 inst_18361 ( .A(net_18208), .Z(net_18209) );
AND4_X4 inst_9032 ( .A2(net_3330), .A1(net_3194), .ZN(net_2663), .A4(net_578), .A3(net_539) );
CLKBUF_X2 inst_14043 ( .A(net_13890), .Z(net_13891) );
OAI21_X2 inst_3065 ( .B2(net_8227), .B1(net_4850), .ZN(net_4735), .A(net_2595) );
SDFF_X2 inst_715 ( .SI(net_8655), .Q(net_8655), .D(net_3954), .SE(net_3885), .CK(net_10061) );
INV_X4 inst_5206 ( .A(net_2467), .ZN(net_2394) );
CLKBUF_X2 inst_14936 ( .A(net_14783), .Z(net_14784) );
CLKBUF_X2 inst_18890 ( .A(net_17190), .Z(net_18738) );
INV_X2 inst_6354 ( .ZN(net_2221), .A(net_2220) );
DFFR_X2 inst_7333 ( .QN(net_7346), .D(net_3258), .CK(net_9555), .RN(x6501) );
AOI21_X2 inst_8941 ( .A(net_5746), .ZN(net_5698), .B2(net_5521), .B1(net_4534) );
INV_X4 inst_5213 ( .ZN(net_2748), .A(net_2220) );
CLKBUF_X2 inst_14113 ( .A(net_11505), .Z(net_13961) );
SDFF_X2 inst_1682 ( .Q(net_8036), .D(net_8036), .SI(net_2710), .SE(net_2545), .CK(net_16473) );
INV_X4 inst_5077 ( .ZN(net_5848), .A(net_5794) );
CLKBUF_X2 inst_18810 ( .A(net_18657), .Z(net_18658) );
CLKBUF_X2 inst_10630 ( .A(net_10477), .Z(net_10478) );
CLKBUF_X2 inst_13778 ( .A(net_13625), .Z(net_13626) );
CLKBUF_X2 inst_18191 ( .A(net_9524), .Z(net_18039) );
NOR2_X2 inst_3505 ( .A1(net_7419), .ZN(net_6220), .A2(net_1766) );
XOR2_X2 inst_31 ( .A(net_6796), .B(net_4373), .Z(net_1208) );
CLKBUF_X2 inst_15136 ( .A(net_14983), .Z(net_14984) );
CLKBUF_X2 inst_15751 ( .A(net_13655), .Z(net_15599) );
CLKBUF_X2 inst_10937 ( .A(net_10467), .Z(net_10785) );
CLKBUF_X2 inst_12730 ( .A(net_12577), .Z(net_12578) );
NOR2_X2 inst_3537 ( .A2(net_2652), .ZN(net_1998), .A1(net_861) );
CLKBUF_X2 inst_9787 ( .A(net_9634), .Z(net_9635) );
CLKBUF_X2 inst_12606 ( .A(net_9253), .Z(net_12454) );
NAND2_X2 inst_4556 ( .A1(net_6385), .A2(net_6184), .ZN(net_3254) );
CLKBUF_X2 inst_19157 ( .A(net_9627), .Z(net_19005) );
CLKBUF_X2 inst_14449 ( .A(net_12668), .Z(net_14297) );
SDFF_X2 inst_1833 ( .D(net_7302), .SI(net_6879), .Q(net_6879), .SE(net_6282), .CK(net_15415) );
SDFFR_X2 inst_2122 ( .SI(net_7184), .Q(net_7184), .D(net_6435), .SE(net_4362), .CK(net_13736), .RN(x6501) );
INV_X4 inst_5301 ( .A(net_1599), .ZN(net_1585) );
AOI22_X2 inst_8160 ( .B1(net_8778), .A1(net_8519), .ZN(net_6240), .A2(net_3861), .B2(net_3860) );
NOR2_X2 inst_3520 ( .ZN(net_1744), .A1(net_1743), .A2(net_1742) );
CLKBUF_X2 inst_9809 ( .A(net_9656), .Z(net_9657) );
CLKBUF_X2 inst_11601 ( .A(net_11448), .Z(net_11449) );
CLKBUF_X2 inst_13041 ( .A(net_12888), .Z(net_12889) );
NOR2_X2 inst_3573 ( .ZN(net_3318), .A1(net_1151), .A2(net_1150) );
CLKBUF_X2 inst_17739 ( .A(net_10795), .Z(net_17587) );
SDFF_X2 inst_623 ( .SI(net_8535), .Q(net_8535), .SE(net_3979), .D(net_3944), .CK(net_10006) );
CLKBUF_X2 inst_11306 ( .A(net_11153), .Z(net_11154) );
CLKBUF_X2 inst_13453 ( .A(net_9130), .Z(net_13301) );
CLKBUF_X2 inst_15612 ( .A(net_15459), .Z(net_15460) );
AOI22_X2 inst_8557 ( .ZN(net_2817), .A1(net_2762), .B2(net_2556), .A2(net_2503), .B1(net_2242) );
SDFF_X2 inst_1621 ( .Q(net_8164), .D(net_8164), .SI(net_2590), .SE(net_2538), .CK(net_15991) );
CLKBUF_X2 inst_10373 ( .A(net_9106), .Z(net_10221) );
CLKBUF_X2 inst_18881 ( .A(net_13049), .Z(net_18729) );
CLKBUF_X2 inst_14877 ( .A(net_10508), .Z(net_14725) );
NOR4_X2 inst_3226 ( .ZN(net_2336), .A4(net_2087), .A3(net_1720), .A2(net_1003), .A1(net_792) );
AOI22_X2 inst_8435 ( .B1(net_6599), .A1(net_6566), .A2(net_6257), .B2(net_6110), .ZN(net_3506) );
CLKBUF_X2 inst_10674 ( .A(net_9939), .Z(net_10522) );
CLKBUF_X2 inst_9609 ( .A(net_9456), .Z(net_9457) );
CLKBUF_X2 inst_13224 ( .A(net_13071), .Z(net_13072) );
CLKBUF_X2 inst_15523 ( .A(net_10590), .Z(net_15371) );
OAI21_X2 inst_3125 ( .B2(net_2299), .ZN(net_2254), .A(net_2253), .B1(net_1133) );
CLKBUF_X2 inst_10571 ( .A(net_10418), .Z(net_10419) );
CLKBUF_X2 inst_14130 ( .A(net_13977), .Z(net_13978) );
CLKBUF_X2 inst_16494 ( .A(net_16341), .Z(net_16342) );
CLKBUF_X2 inst_18998 ( .A(net_18845), .Z(net_18846) );
CLKBUF_X2 inst_16546 ( .A(net_16393), .Z(net_16394) );
SDFF_X2 inst_760 ( .Q(net_8802), .D(net_8802), .SI(net_3955), .SE(net_3879), .CK(net_10985) );
CLKBUF_X2 inst_10562 ( .A(net_10409), .Z(net_10410) );
CLKBUF_X2 inst_10750 ( .A(net_10597), .Z(net_10598) );
CLKBUF_X2 inst_10814 ( .A(net_10661), .Z(net_10662) );
CLKBUF_X2 inst_12842 ( .A(net_12689), .Z(net_12690) );
AOI21_X4 inst_8867 ( .B1(net_6147), .ZN(net_4506), .B2(net_4403), .A(net_4358) );
CLKBUF_X2 inst_18799 ( .A(net_18646), .Z(net_18647) );
SDFF_X2 inst_1696 ( .Q(net_8162), .D(net_8162), .SI(net_2575), .SE(net_2538), .CK(net_15974) );
CLKBUF_X2 inst_15863 ( .A(net_12811), .Z(net_15711) );
CLKBUF_X2 inst_16591 ( .A(net_16438), .Z(net_16439) );
CLKBUF_X2 inst_14519 ( .A(net_9989), .Z(net_14367) );
CLKBUF_X2 inst_9347 ( .A(net_9194), .Z(net_9195) );
CLKBUF_X2 inst_17171 ( .A(net_17018), .Z(net_17019) );
CLKBUF_X2 inst_17203 ( .A(net_13172), .Z(net_17051) );
NAND4_X2 inst_3727 ( .ZN(net_4303), .A1(net_4154), .A2(net_4153), .A3(net_4152), .A4(net_4151) );
CLKBUF_X2 inst_9831 ( .A(net_9302), .Z(net_9679) );
CLKBUF_X2 inst_10812 ( .A(net_10659), .Z(net_10660) );
CLKBUF_X2 inst_12237 ( .A(net_12084), .Z(net_12085) );
CLKBUF_X2 inst_17189 ( .A(net_17036), .Z(net_17037) );
DFFR_X2 inst_7258 ( .QN(net_7308), .D(net_1997), .CK(net_15933), .RN(x6501) );
NAND3_X2 inst_3989 ( .A2(net_9048), .ZN(net_3976), .A1(net_1593), .A3(net_1592) );
CLKBUF_X2 inst_10000 ( .A(net_9847), .Z(net_9848) );
CLKBUF_X2 inst_14973 ( .A(net_14376), .Z(net_14821) );
CLKBUF_X2 inst_12934 ( .A(net_12781), .Z(net_12782) );
NOR2_X2 inst_3569 ( .A1(net_7519), .ZN(net_1527), .A2(net_832) );
DFFR_X2 inst_7268 ( .QN(net_7405), .D(net_1980), .CK(net_17855), .RN(x6501) );
NOR2_X2 inst_3411 ( .ZN(net_3374), .A1(net_3259), .A2(net_3220) );
CLKBUF_X2 inst_10436 ( .A(net_10283), .Z(net_10284) );
SDFFR_X2 inst_2524 ( .D(net_7373), .SE(net_2387), .SI(net_288), .Q(net_288), .CK(net_16388), .RN(x6501) );
SDFF_X2 inst_1446 ( .SI(net_7294), .Q(net_7111), .D(net_7111), .SE(net_6278), .CK(net_17708) );
CLKBUF_X2 inst_9486 ( .A(net_9333), .Z(net_9334) );
SDFFR_X2 inst_2421 ( .SE(net_2683), .D(net_2681), .SI(net_468), .Q(net_468), .CK(net_13939), .RN(x6501) );
SDFF_X2 inst_390 ( .Q(net_8837), .D(net_8837), .SE(net_3964), .SI(net_3963), .CK(net_10945) );
CLKBUF_X2 inst_16866 ( .A(net_11303), .Z(net_16714) );
CLKBUF_X2 inst_17754 ( .A(net_17601), .Z(net_17602) );
SDFF_X2 inst_1062 ( .D(net_7322), .SI(net_6630), .Q(net_6630), .SE(net_3123), .CK(net_9153) );
AOI22_X2 inst_8181 ( .B1(net_8827), .A1(net_8346), .A2(net_6265), .B2(net_6253), .ZN(net_3851) );
CLKBUF_X2 inst_14455 ( .A(net_14302), .Z(net_14303) );
CLKBUF_X2 inst_16669 ( .A(net_14604), .Z(net_16517) );
AOI22_X2 inst_7996 ( .A1(net_7961), .B1(net_7791), .A2(net_6092), .B2(net_6091), .ZN(net_4137) );
CLKBUF_X2 inst_13757 ( .A(net_12239), .Z(net_13605) );
CLKBUF_X2 inst_12814 ( .A(net_10321), .Z(net_12662) );
CLKBUF_X2 inst_14361 ( .A(net_14208), .Z(net_14209) );
CLKBUF_X2 inst_16745 ( .A(net_16592), .Z(net_16593) );
CLKBUF_X2 inst_10277 ( .A(net_10124), .Z(net_10125) );
CLKBUF_X2 inst_15944 ( .A(net_12618), .Z(net_15792) );
CLKBUF_X2 inst_12440 ( .A(net_12287), .Z(net_12288) );
DFFR_X2 inst_7063 ( .QN(net_7193), .D(net_4312), .CK(net_13737), .RN(x6501) );
SDFFR_X1 inst_2642 ( .D(net_6765), .SE(net_4506), .CK(net_9254), .RN(x6501), .SI(x1912), .Q(x1912) );
CLKBUF_X2 inst_12539 ( .A(net_10400), .Z(net_12387) );
CLKBUF_X2 inst_15974 ( .A(net_15821), .Z(net_15822) );
CLKBUF_X2 inst_18817 ( .A(net_12967), .Z(net_18665) );
CLKBUF_X2 inst_18317 ( .A(net_18164), .Z(net_18165) );
CLKBUF_X2 inst_18995 ( .A(net_18842), .Z(net_18843) );
CLKBUF_X2 inst_14394 ( .A(net_14241), .Z(net_14242) );
XNOR2_X2 inst_123 ( .ZN(net_2929), .A(net_2808), .B(net_847) );
INV_X4 inst_5250 ( .A(net_2129), .ZN(net_1858) );
SDFFR_X2 inst_2160 ( .QN(net_7577), .D(net_3944), .SE(net_3144), .SI(net_529), .CK(net_10877), .RN(x6501) );
INV_X4 inst_5181 ( .ZN(net_2869), .A(net_2817) );
CLKBUF_X2 inst_10981 ( .A(net_10828), .Z(net_10829) );
SDFFR_X2 inst_2298 ( .D(net_4459), .SE(net_2757), .SI(net_419), .Q(net_419), .CK(net_17296), .RN(x6501) );
CLKBUF_X2 inst_14355 ( .A(net_14202), .Z(net_14203) );
CLKBUF_X2 inst_14546 ( .A(net_14393), .Z(net_14394) );
XNOR2_X2 inst_167 ( .ZN(net_1826), .A(net_1594), .B(net_1539) );
CLKBUF_X2 inst_11660 ( .A(net_11507), .Z(net_11508) );
CLKBUF_X2 inst_11354 ( .A(net_11201), .Z(net_11202) );
CLKBUF_X2 inst_13138 ( .A(net_12985), .Z(net_12986) );
NAND2_X1 inst_4913 ( .A1(net_6807), .A2(net_6804), .ZN(net_605) );
AOI22_X2 inst_8524 ( .B1(net_6523), .A1(net_6490), .A2(net_6137), .B2(net_6104), .ZN(net_3416) );
SDFFR_X2 inst_2475 ( .Q(net_8981), .D(net_8981), .SI(net_2594), .SE(net_2562), .CK(net_13925), .RN(x6501) );
NAND2_X2 inst_4874 ( .ZN(net_1070), .A1(x2805), .A2(x2746) );
DFF_X1 inst_6824 ( .Q(net_8219), .D(net_4443), .CK(net_17197) );
CLKBUF_X2 inst_13033 ( .A(net_12571), .Z(net_12881) );
CLKBUF_X2 inst_17848 ( .A(net_17695), .Z(net_17696) );
AND2_X2 inst_9195 ( .ZN(net_1569), .A1(net_1568), .A2(net_1567) );
CLKBUF_X2 inst_13131 ( .A(net_12978), .Z(net_12979) );
XNOR2_X2 inst_331 ( .B(net_7388), .A(net_6370), .ZN(net_812) );
CLKBUF_X2 inst_10691 ( .A(net_9642), .Z(net_10539) );
CLKBUF_X2 inst_13312 ( .A(net_11598), .Z(net_13160) );
AOI21_X2 inst_8948 ( .A(net_5783), .ZN(net_5675), .B1(net_5472), .B2(net_5266) );
CLKBUF_X2 inst_14317 ( .A(net_9118), .Z(net_14165) );
CLKBUF_X2 inst_11227 ( .A(net_11074), .Z(net_11075) );
SDFFR_X2 inst_2353 ( .D(net_2728), .SE(net_2313), .SI(net_447), .Q(net_447), .CK(net_16542), .RN(x6501) );
CLKBUF_X2 inst_11921 ( .A(net_9751), .Z(net_11769) );
CLKBUF_X2 inst_17552 ( .A(net_14305), .Z(net_17400) );
CLKBUF_X2 inst_13483 ( .A(net_9519), .Z(net_13331) );
SDFFR_X1 inst_2762 ( .QN(net_9010), .D(net_6165), .SE(net_3144), .SI(net_2246), .CK(net_11128), .RN(x6501) );
SDFF_X2 inst_997 ( .D(net_7336), .SI(net_6644), .Q(net_6644), .SE(net_3123), .CK(net_9499) );
SDFF_X2 inst_857 ( .SI(net_8637), .Q(net_8637), .D(net_3981), .SE(net_3885), .CK(net_12941) );
CLKBUF_X2 inst_16235 ( .A(net_13809), .Z(net_16083) );
NAND2_X2 inst_4824 ( .A2(net_7401), .ZN(net_1369), .A1(net_669) );
INV_X2 inst_6403 ( .A(net_2530), .ZN(net_1128) );
NAND2_X2 inst_4179 ( .ZN(net_5325), .A1(net_5077), .A2(net_5076) );
CLKBUF_X2 inst_12721 ( .A(net_10140), .Z(net_12569) );
INV_X4 inst_5951 ( .A(net_6349), .ZN(net_970) );
NAND3_X2 inst_4006 ( .A3(net_1536), .A2(net_1515), .ZN(net_1261), .A1(net_906) );
AOI22_X2 inst_7988 ( .A1(net_7960), .B1(net_7790), .A2(net_6092), .B2(net_6091), .ZN(net_4144) );
CLKBUF_X2 inst_15918 ( .A(net_15765), .Z(net_15766) );
CLKBUF_X2 inst_18532 ( .A(net_18379), .Z(net_18380) );
OAI211_X2 inst_3203 ( .B(net_5955), .C2(net_2876), .ZN(net_2420), .A(net_912), .C1(net_911) );
CLKBUF_X2 inst_15368 ( .A(net_15215), .Z(net_15216) );
INV_X4 inst_5073 ( .ZN(net_5855), .A(net_5808) );
CLKBUF_X2 inst_13951 ( .A(net_10883), .Z(net_13799) );
SDFF_X2 inst_1310 ( .Q(net_8090), .D(net_8090), .SE(net_2707), .SI(net_2574), .CK(net_16079) );
NOR3_X2 inst_3280 ( .ZN(net_2794), .A1(net_2400), .A3(net_2396), .A2(net_1494) );
NAND2_X2 inst_4491 ( .A1(net_7203), .A2(net_5655), .ZN(net_4481) );
DFFR_X1 inst_7397 ( .D(net_5828), .CK(net_17171), .RN(x6501), .Q(x170) );
OR2_X4 inst_2823 ( .A2(net_6206), .ZN(net_4406), .A1(net_4320) );
CLKBUF_X2 inst_11594 ( .A(net_10067), .Z(net_11442) );
CLKBUF_X2 inst_13981 ( .A(net_13828), .Z(net_13829) );
CLKBUF_X2 inst_13413 ( .A(net_12396), .Z(net_13261) );
CLKBUF_X2 inst_15171 ( .A(net_15018), .Z(net_15019) );
CLKBUF_X2 inst_16711 ( .A(net_16558), .Z(net_16559) );
CLKBUF_X2 inst_14464 ( .A(net_14311), .Z(net_14312) );
XNOR2_X2 inst_136 ( .ZN(net_2745), .A(net_2553), .B(net_2549) );
INV_X4 inst_5839 ( .A(net_8963), .ZN(net_1061) );
CLKBUF_X2 inst_11733 ( .A(net_9621), .Z(net_11581) );
CLKBUF_X2 inst_13837 ( .A(net_10835), .Z(net_13685) );
SDFF_X2 inst_1526 ( .Q(net_7900), .D(net_7900), .SI(net_2710), .SE(net_2543), .CK(net_16508) );
SDFFR_X2 inst_2547 ( .QN(net_6348), .SE(net_2147), .D(net_2137), .SI(net_1615), .CK(net_18325), .RN(x6501) );
NAND2_X2 inst_4637 ( .A2(net_6264), .ZN(net_6218), .A1(net_5691) );
CLKBUF_X2 inst_16800 ( .A(net_16647), .Z(net_16648) );
SDFF_X2 inst_1047 ( .SI(net_7311), .Q(net_6685), .D(net_6685), .SE(net_3125), .CK(net_12105) );
CLKBUF_X2 inst_15790 ( .A(net_15637), .Z(net_15638) );
DFFS_X2 inst_6860 ( .QN(net_7351), .D(net_5527), .CK(net_9548), .SN(x6501) );
AOI22_X2 inst_8507 ( .B1(net_6588), .A1(net_6555), .A2(net_6257), .B2(net_6110), .ZN(net_3433) );
CLKBUF_X2 inst_11768 ( .A(net_11615), .Z(net_11616) );
NAND4_X2 inst_3700 ( .ZN(net_4437), .A4(net_4339), .A1(net_3764), .A2(net_3763), .A3(net_3762) );
DFF_X1 inst_6744 ( .QN(net_6788), .D(net_5625), .CK(net_11583) );
CLKBUF_X2 inst_12432 ( .A(net_12279), .Z(net_12280) );
CLKBUF_X2 inst_15519 ( .A(net_15189), .Z(net_15367) );
CLKBUF_X2 inst_16955 ( .A(net_12766), .Z(net_16803) );
SDFF_X2 inst_1858 ( .D(net_7286), .SI(net_6943), .Q(net_6943), .SE(net_6281), .CK(net_17678) );
CLKBUF_X2 inst_17120 ( .A(net_16967), .Z(net_16968) );
NAND4_X2 inst_3846 ( .A4(net_7223), .ZN(net_2400), .A2(net_2085), .A1(net_1802), .A3(net_769) );
CLKBUF_X2 inst_13668 ( .A(net_13515), .Z(net_13516) );
SDFF_X2 inst_1334 ( .SI(net_7683), .Q(net_7683), .D(net_2720), .SE(net_2714), .CK(net_18081) );
CLKBUF_X2 inst_17491 ( .A(net_17338), .Z(net_17339) );
INV_X4 inst_5944 ( .A(net_7303), .ZN(net_827) );
INV_X4 inst_5383 ( .A(net_1431), .ZN(net_1105) );
INV_X4 inst_6129 ( .A(net_7508), .ZN(net_3334) );
CLKBUF_X2 inst_14735 ( .A(net_14582), .Z(net_14583) );
DFFR_X2 inst_7273 ( .QN(net_6392), .D(net_2035), .CK(net_15669), .RN(x6501) );
CLKBUF_X2 inst_12130 ( .A(net_11691), .Z(net_11978) );
CLKBUF_X2 inst_15567 ( .A(net_15414), .Z(net_15415) );
CLKBUF_X2 inst_11453 ( .A(net_10252), .Z(net_11301) );
XNOR2_X2 inst_265 ( .A(net_7581), .B(net_3581), .ZN(net_1115) );
SDFF_X2 inst_2055 ( .SI(net_7803), .Q(net_7803), .D(net_2716), .SE(net_2459), .CK(net_17042) );
CLKBUF_X2 inst_11702 ( .A(net_10056), .Z(net_11550) );
AOI22_X2 inst_7783 ( .A1(net_5268), .B2(net_5267), .ZN(net_4868), .A2(net_4632), .B1(net_182) );
INV_X4 inst_5554 ( .ZN(net_831), .A(net_635) );
CLKBUF_X2 inst_18667 ( .A(net_10983), .Z(net_18515) );
NOR3_X2 inst_3262 ( .ZN(net_3212), .A1(net_3148), .A3(net_2020), .A2(net_1742) );
CLKBUF_X2 inst_17932 ( .A(net_17779), .Z(net_17780) );
NAND2_X2 inst_4566 ( .ZN(net_3220), .A1(net_3030), .A2(net_2994) );
CLKBUF_X2 inst_12993 ( .A(net_12840), .Z(net_12841) );
CLKBUF_X2 inst_10653 ( .A(net_10500), .Z(net_10501) );
INV_X2 inst_6301 ( .ZN(net_3992), .A(net_3906) );
DFFR_X2 inst_7249 ( .QN(net_7259), .D(net_2061), .CK(net_15051), .RN(x6501) );
AOI22_X2 inst_7975 ( .A1(net_7958), .B1(net_7788), .A2(net_6092), .B2(net_6091), .ZN(net_4155) );
NAND3_X2 inst_3954 ( .ZN(net_3217), .A2(net_3072), .A1(net_3002), .A3(net_2990) );
CLKBUF_X2 inst_12956 ( .A(net_11628), .Z(net_12804) );
CLKBUF_X2 inst_9367 ( .A(net_9214), .Z(net_9215) );
XNOR2_X2 inst_222 ( .ZN(net_1390), .A(net_1389), .B(net_648) );
CLKBUF_X2 inst_18857 ( .A(net_18704), .Z(net_18705) );
INV_X2 inst_6372 ( .A(net_1733), .ZN(net_1627) );
INV_X4 inst_6073 ( .A(net_7490), .ZN(net_4697) );
CLKBUF_X2 inst_13166 ( .A(net_13013), .Z(net_13014) );
CLKBUF_X2 inst_12218 ( .A(net_9599), .Z(net_12066) );
DFF_X1 inst_6728 ( .Q(net_6774), .D(net_5641), .CK(net_9216) );
SDFF_X2 inst_1302 ( .Q(net_7820), .D(net_7820), .SE(net_2730), .SI(net_2589), .CK(net_15629) );
CLKBUF_X2 inst_18220 ( .A(net_16296), .Z(net_18068) );
CLKBUF_X2 inst_10609 ( .A(net_10456), .Z(net_10457) );
SDFF_X2 inst_1648 ( .SI(net_7728), .Q(net_7728), .D(net_2717), .SE(net_2559), .CK(net_16477) );
SDFF_X2 inst_1079 ( .D(net_7312), .SI(net_6488), .Q(net_6488), .SE(net_3071), .CK(net_12010) );
INV_X4 inst_5847 ( .A(net_6378), .ZN(net_948) );
CLKBUF_X2 inst_13958 ( .A(net_13805), .Z(net_13806) );
CLKBUF_X2 inst_13833 ( .A(net_12176), .Z(net_13681) );
CLKBUF_X2 inst_19144 ( .A(net_17753), .Z(net_18992) );
CLKBUF_X2 inst_16857 ( .A(net_16704), .Z(net_16705) );
NAND3_X2 inst_3925 ( .ZN(net_5613), .A1(net_5542), .A3(net_5476), .A2(net_5291) );
CLKBUF_X2 inst_18918 ( .A(net_18765), .Z(net_18766) );
SDFFR_X2 inst_2606 ( .D(net_7374), .Q(net_7271), .SI(net_1808), .SE(net_1327), .CK(net_17508), .RN(x6501) );
NAND2_X2 inst_4314 ( .A1(net_7137), .A2(net_5166), .ZN(net_5143) );
CLKBUF_X2 inst_9837 ( .A(net_9149), .Z(net_9685) );
SDFFR_X2 inst_2523 ( .D(net_7370), .SE(net_2387), .SI(net_285), .Q(net_285), .CK(net_16391), .RN(x6501) );
SDFF_X2 inst_506 ( .SI(net_8600), .Q(net_8600), .SE(net_3984), .D(net_3981), .CK(net_12996) );
CLKBUF_X2 inst_10662 ( .A(net_10509), .Z(net_10510) );
CLKBUF_X2 inst_13569 ( .A(net_13416), .Z(net_13417) );
CLKBUF_X2 inst_17834 ( .A(net_17681), .Z(net_17682) );
CLKBUF_X2 inst_11782 ( .A(net_11606), .Z(net_11630) );
AOI22_X2 inst_8572 ( .B1(net_2800), .A1(net_2701), .ZN(net_1920), .A2(net_1919), .B2(net_1918) );
CLKBUF_X2 inst_10835 ( .A(net_10682), .Z(net_10683) );
SDFF_X2 inst_1323 ( .Q(net_7807), .D(net_7807), .SE(net_2730), .SI(net_2585), .CK(net_15852) );
SDFF_X2 inst_1085 ( .D(net_7339), .SI(net_6515), .Q(net_6515), .SE(net_3071), .CK(net_11888) );
CLKBUF_X2 inst_14048 ( .A(net_10330), .Z(net_13896) );
CLKBUF_X2 inst_18177 ( .A(net_13287), .Z(net_18025) );
AOI221_X2 inst_8791 ( .C1(net_7201), .C2(net_5655), .B2(net_4965), .ZN(net_4910), .A(net_4908), .B1(net_303) );
CLKBUF_X2 inst_10464 ( .A(net_10311), .Z(net_10312) );
SDFFR_X1 inst_2655 ( .D(net_6777), .SE(net_4506), .CK(net_9232), .RN(x6501), .SI(x1575), .Q(x1575) );
SDFF_X2 inst_1720 ( .Q(net_8007), .D(net_8007), .SI(net_2716), .SE(net_2542), .CK(net_16822) );
XNOR2_X2 inst_160 ( .ZN(net_1850), .B(net_1760), .A(net_1759) );
AOI21_X2 inst_8889 ( .B2(net_5871), .ZN(net_5808), .A(net_5807), .B1(net_2671) );
CLKBUF_X2 inst_14420 ( .A(net_14267), .Z(net_14268) );
CLKBUF_X2 inst_9243 ( .A(net_9062), .Z(net_9091) );
CLKBUF_X2 inst_18494 ( .A(net_15005), .Z(net_18342) );
SDFF_X2 inst_370 ( .SI(net_8541), .Q(net_8541), .SE(net_3979), .D(net_3963), .CK(net_12367) );
DFFR_X1 inst_7450 ( .QN(net_8933), .D(net_4749), .CK(net_17310), .RN(x6501) );
AOI22_X2 inst_7825 ( .A2(net_5535), .B2(net_5260), .ZN(net_4698), .B1(net_4697), .A1(net_449) );
CLKBUF_X2 inst_10414 ( .A(net_10261), .Z(net_10262) );
SDFF_X2 inst_1265 ( .Q(net_8111), .D(net_8111), .SE(net_2707), .SI(net_2703), .CK(net_14032) );
CLKBUF_X2 inst_14480 ( .A(net_11906), .Z(net_14328) );
CLKBUF_X2 inst_10669 ( .A(net_10088), .Z(net_10517) );
AOI22_X2 inst_8371 ( .B1(net_8781), .A1(net_8522), .A2(net_3861), .B2(net_3860), .ZN(net_3677) );
AOI22_X2 inst_8176 ( .B1(net_8678), .A1(net_8641), .B2(net_6109), .A2(net_3857), .ZN(net_3854) );
CLKBUF_X2 inst_11288 ( .A(net_11135), .Z(net_11136) );
SDFF_X2 inst_1321 ( .SI(net_7693), .Q(net_7693), .D(net_2749), .SE(net_2714), .CK(net_14436) );
SDFF_X2 inst_1012 ( .SI(net_7326), .Q(net_6667), .D(net_6667), .SE(net_3126), .CK(net_11296) );
INV_X4 inst_5255 ( .ZN(net_2066), .A(net_1880) );
CLKBUF_X2 inst_12768 ( .A(net_12615), .Z(net_12616) );
CLKBUF_X2 inst_16082 ( .A(net_15929), .Z(net_15930) );
AOI22_X2 inst_8341 ( .A1(net_8626), .B1(net_8441), .A2(net_3864), .B2(net_3863), .ZN(net_3706) );
NOR2_X2 inst_3492 ( .A1(net_2074), .ZN(net_2067), .A2(net_2066) );
CLKBUF_X2 inst_18542 ( .A(net_18389), .Z(net_18390) );
CLKBUF_X2 inst_14032 ( .A(net_13879), .Z(net_13880) );
CLKBUF_X2 inst_14724 ( .A(net_14571), .Z(net_14572) );
AOI211_X2 inst_9015 ( .ZN(net_2202), .B(net_1911), .C2(net_1740), .A(net_1664), .C1(net_1595) );
OAI21_X2 inst_3149 ( .B2(net_2048), .ZN(net_1987), .A(net_1972), .B1(net_649) );
CLKBUF_X2 inst_17644 ( .A(net_17491), .Z(net_17492) );
NAND2_X4 inst_4034 ( .A2(net_6157), .A1(net_6100), .ZN(net_2911) );
SDFF_X2 inst_377 ( .SI(net_8380), .Q(net_8380), .SE(net_3969), .D(net_3946), .CK(net_10774) );
CLKBUF_X2 inst_13570 ( .A(net_13417), .Z(net_13418) );
DFFR_X2 inst_6993 ( .QN(net_6312), .D(net_5849), .CK(net_16950), .RN(x6501) );
CLKBUF_X2 inst_10157 ( .A(net_10004), .Z(net_10005) );
NAND3_X2 inst_3946 ( .ZN(net_4379), .A3(net_4324), .A2(net_4322), .A1(net_4317) );
NAND2_X2 inst_4760 ( .ZN(net_2435), .A1(net_394), .A2(net_391) );
CLKBUF_X2 inst_15703 ( .A(net_15550), .Z(net_15551) );
NAND3_X2 inst_3920 ( .ZN(net_5618), .A1(net_5547), .A3(net_5481), .A2(net_5311) );
DFFS_X1 inst_6953 ( .D(net_3231), .CK(net_16337), .SN(x6501), .Q(x898) );
DFFS_X1 inst_6920 ( .D(net_6145), .CK(net_13666), .SN(x6501), .Q(x778) );
OAI21_X2 inst_3018 ( .B2(net_5044), .ZN(net_5042), .A(net_4887), .B1(net_1676) );
OAI21_X2 inst_3078 ( .ZN(net_4222), .A(net_3548), .B2(net_3245), .B1(net_1111) );
CLKBUF_X2 inst_13750 ( .A(net_13597), .Z(net_13598) );
INV_X4 inst_5792 ( .A(net_9009), .ZN(net_546) );
CLKBUF_X2 inst_12779 ( .A(net_12626), .Z(net_12627) );
CLKBUF_X2 inst_9731 ( .A(net_9100), .Z(net_9579) );
CLKBUF_X2 inst_13579 ( .A(net_13426), .Z(net_13427) );
CLKBUF_X2 inst_18481 ( .A(net_18328), .Z(net_18329) );
INV_X8 inst_5054 ( .A(net_6261), .ZN(net_6259) );
INV_X4 inst_5926 ( .ZN(net_2741), .A(net_278) );
CLKBUF_X2 inst_16113 ( .A(net_15960), .Z(net_15961) );
NAND2_X2 inst_4627 ( .ZN(net_2775), .A1(net_2529), .A2(net_2444) );
CLKBUF_X2 inst_17018 ( .A(net_16865), .Z(net_16866) );
CLKBUF_X2 inst_12414 ( .A(net_12261), .Z(net_12262) );
CLKBUF_X2 inst_13559 ( .A(net_13406), .Z(net_13407) );
CLKBUF_X2 inst_14429 ( .A(net_14276), .Z(net_14277) );
CLKBUF_X2 inst_16110 ( .A(net_15957), .Z(net_15958) );
XNOR2_X2 inst_107 ( .ZN(net_5712), .A(net_5467), .B(net_2289) );
CLKBUF_X2 inst_14191 ( .A(net_9737), .Z(net_14039) );
CLKBUF_X2 inst_16166 ( .A(net_13723), .Z(net_16014) );
SDFF_X2 inst_990 ( .D(net_7328), .SI(net_6636), .Q(net_6636), .SE(net_3123), .CK(net_9528) );
CLKBUF_X2 inst_12381 ( .A(net_12228), .Z(net_12229) );
CLKBUF_X2 inst_16807 ( .A(net_16654), .Z(net_16655) );
DFFR_X2 inst_7225 ( .QN(net_8967), .D(net_2238), .CK(net_16293), .RN(x6501) );
CLKBUF_X2 inst_10412 ( .A(net_10259), .Z(net_10260) );
NAND2_X2 inst_4710 ( .A2(net_6408), .ZN(net_2217), .A1(net_1843) );
NAND4_X2 inst_3628 ( .ZN(net_5590), .A2(net_5459), .A1(net_5283), .A4(net_4777), .A3(net_4502) );
CLKBUF_X2 inst_15632 ( .A(net_15479), .Z(net_15480) );
SDFFR_X2 inst_2366 ( .SE(net_2260), .Q(net_331), .D(net_331), .CK(net_9300), .RN(x6501), .SI(x2594) );
CLKBUF_X2 inst_10093 ( .A(net_9940), .Z(net_9941) );
CLKBUF_X2 inst_14886 ( .A(net_14262), .Z(net_14734) );
INV_X8 inst_5049 ( .ZN(net_6275), .A(net_6190) );
CLKBUF_X2 inst_11343 ( .A(net_10890), .Z(net_11191) );
CLKBUF_X2 inst_14155 ( .A(net_14002), .Z(net_14003) );
CLKBUF_X2 inst_13998 ( .A(net_12047), .Z(net_13846) );
NAND2_X2 inst_4605 ( .A2(net_6144), .ZN(net_2631), .A1(net_2630) );
CLKBUF_X2 inst_10351 ( .A(net_10198), .Z(net_10199) );
CLKBUF_X2 inst_11207 ( .A(net_11054), .Z(net_11055) );
SDFF_X2 inst_1237 ( .Q(net_7953), .D(net_7953), .SE(net_2755), .SI(net_2706), .CK(net_18899) );
CLKBUF_X2 inst_12873 ( .A(net_12475), .Z(net_12721) );
CLKBUF_X2 inst_15196 ( .A(net_11812), .Z(net_15044) );
DFFR_X2 inst_7175 ( .D(net_2523), .QN(net_401), .CK(net_14828), .RN(x6501) );
NOR3_X2 inst_3310 ( .ZN(net_1743), .A1(net_1222), .A3(net_994), .A2(net_964) );
OAI21_X2 inst_3062 ( .B2(net_8248), .B1(net_4850), .ZN(net_4742), .A(net_2629) );
INV_X2 inst_6267 ( .A(net_8249), .ZN(net_4630) );
CLKBUF_X2 inst_14249 ( .A(net_14096), .Z(net_14097) );
CLKBUF_X2 inst_13459 ( .A(net_13306), .Z(net_13307) );
INV_X4 inst_5100 ( .ZN(net_5693), .A(net_5663) );
AOI22_X2 inst_8536 ( .B1(net_6526), .A1(net_6493), .A2(net_6137), .B2(net_6104), .ZN(net_3404) );
CLKBUF_X2 inst_15239 ( .A(net_15086), .Z(net_15087) );
CLKBUF_X2 inst_13967 ( .A(net_13814), .Z(net_13815) );
CLKBUF_X2 inst_14745 ( .A(net_14592), .Z(net_14593) );
INV_X4 inst_6013 ( .A(net_7416), .ZN(net_1444) );
SDFF_X2 inst_383 ( .SI(net_8388), .Q(net_8388), .SE(net_3969), .D(net_3967), .CK(net_13070) );
CLKBUF_X2 inst_15017 ( .A(net_14864), .Z(net_14865) );
CLKBUF_X2 inst_11793 ( .A(net_11640), .Z(net_11641) );
CLKBUF_X2 inst_13561 ( .A(net_13408), .Z(net_13409) );
NAND2_X2 inst_4132 ( .ZN(net_5391), .A2(net_5222), .A1(net_5123) );
DFFR_X2 inst_7031 ( .QN(net_7489), .D(net_5045), .CK(net_16598), .RN(x6501) );
CLKBUF_X2 inst_9765 ( .A(net_9612), .Z(net_9613) );
CLKBUF_X2 inst_17908 ( .A(net_17755), .Z(net_17756) );
CLKBUF_X2 inst_19115 ( .A(net_18962), .Z(net_18963) );
CLKBUF_X2 inst_16651 ( .A(net_16498), .Z(net_16499) );
CLKBUF_X2 inst_11801 ( .A(net_11648), .Z(net_11649) );
CLKBUF_X2 inst_15972 ( .A(net_15819), .Z(net_15820) );
INV_X4 inst_5372 ( .ZN(net_1343), .A(net_1127) );
NOR2_X2 inst_3375 ( .ZN(net_5550), .A1(net_5325), .A2(net_5324) );
XNOR2_X2 inst_234 ( .A(net_6383), .ZN(net_1250), .B(net_801) );
CLKBUF_X2 inst_16428 ( .A(net_16275), .Z(net_16276) );
INV_X4 inst_5293 ( .ZN(net_1861), .A(net_1309) );
CLKBUF_X2 inst_16893 ( .A(net_16740), .Z(net_16741) );
CLKBUF_X2 inst_12398 ( .A(net_12245), .Z(net_12246) );
CLKBUF_X2 inst_18604 ( .A(net_18451), .Z(net_18452) );
CLKBUF_X2 inst_13975 ( .A(net_11492), .Z(net_13823) );
NOR2_X2 inst_3429 ( .A2(net_5981), .ZN(net_3182), .A1(net_3181) );
SDFF_X2 inst_1328 ( .SI(net_7689), .Q(net_7689), .D(net_2722), .SE(net_2714), .CK(net_14937) );
CLKBUF_X2 inst_18204 ( .A(net_18051), .Z(net_18052) );
AOI22_X2 inst_8429 ( .B1(net_6730), .A1(net_6697), .B2(net_6202), .A2(net_3520), .ZN(net_3512) );
CLKBUF_X2 inst_15434 ( .A(net_11340), .Z(net_15282) );
SDFF_X2 inst_1776 ( .D(net_7276), .SI(net_6853), .Q(net_6853), .SE(net_6282), .CK(net_17383) );
SDFFR_X2 inst_2335 ( .D(net_7368), .SE(net_2738), .SI(net_264), .Q(net_264), .CK(net_13552), .RN(x6501) );
CLKBUF_X2 inst_13157 ( .A(net_11121), .Z(net_13005) );
CLKBUF_X2 inst_18699 ( .A(net_16435), .Z(net_18547) );
SDFF_X2 inst_598 ( .SI(net_8372), .Q(net_8372), .SE(net_3969), .D(net_3943), .CK(net_13125) );
SDFF_X2 inst_1624 ( .Q(net_8167), .D(net_8167), .SI(net_2713), .SE(net_2538), .CK(net_13776) );
CLKBUF_X2 inst_14868 ( .A(net_14715), .Z(net_14716) );
CLKBUF_X2 inst_10595 ( .A(net_10442), .Z(net_10443) );
CLKBUF_X2 inst_10728 ( .A(net_10575), .Z(net_10576) );
OAI21_X2 inst_3167 ( .B1(net_7262), .ZN(net_1996), .A(net_1534), .B2(net_898) );
CLKBUF_X2 inst_13501 ( .A(net_13348), .Z(net_13349) );
CLKBUF_X2 inst_14029 ( .A(net_13876), .Z(net_13877) );
DFFR_X2 inst_7205 ( .D(net_2377), .QN(net_208), .CK(net_17887), .RN(x6501) );
XNOR2_X2 inst_325 ( .B(net_7387), .ZN(net_934), .A(net_933) );
CLKBUF_X2 inst_14861 ( .A(net_14708), .Z(net_14709) );
INV_X2 inst_6502 ( .A(net_5946), .ZN(x1215) );
CLKBUF_X2 inst_16579 ( .A(net_10091), .Z(net_16427) );
AOI221_X2 inst_8858 ( .B1(net_8859), .C1(net_8304), .B2(net_6252), .ZN(net_6235), .C2(net_4345), .A(net_4233) );
NAND2_X2 inst_4769 ( .ZN(net_1837), .A2(net_1670), .A1(x5001) );
SDFF_X2 inst_1197 ( .SI(net_7300), .Q(net_7077), .D(net_7077), .SE(net_6280), .CK(net_18221) );
CLKBUF_X2 inst_18371 ( .A(net_18218), .Z(net_18219) );
DFFS_X1 inst_6958 ( .D(net_2586), .CK(net_16574), .SN(x6501), .Q(x683) );
CLKBUF_X2 inst_10544 ( .A(net_10391), .Z(net_10392) );
SDFF_X2 inst_955 ( .SI(net_7341), .Q(net_6715), .D(net_6715), .SE(net_3125), .CK(net_11920) );
CLKBUF_X2 inst_15793 ( .A(net_15640), .Z(net_15641) );
CLKBUF_X2 inst_11041 ( .A(net_9941), .Z(net_10889) );
CLKBUF_X2 inst_9519 ( .A(net_9165), .Z(net_9367) );
CLKBUF_X2 inst_18264 ( .A(net_18111), .Z(net_18112) );
CLKBUF_X2 inst_15157 ( .A(net_15004), .Z(net_15005) );
INV_X4 inst_5851 ( .A(net_7576), .ZN(net_536) );
CLKBUF_X2 inst_18418 ( .A(net_18265), .Z(net_18266) );
CLKBUF_X2 inst_16364 ( .A(net_11228), .Z(net_16212) );
HA_X1 inst_6665 ( .S(net_3271), .CO(net_3270), .A(net_3269), .B(net_3099) );
CLKBUF_X2 inst_12502 ( .A(net_12349), .Z(net_12350) );
DFFR_X2 inst_7117 ( .QN(net_7614), .D(net_3050), .CK(net_9802), .RN(x6501) );
OR2_X4 inst_2842 ( .A2(net_6094), .ZN(net_2172), .A1(net_844) );
CLKBUF_X2 inst_11142 ( .A(net_10989), .Z(net_10990) );
CLKBUF_X2 inst_13663 ( .A(net_12583), .Z(net_13511) );
NAND4_X2 inst_3792 ( .ZN(net_3634), .A1(net_3521), .A2(net_3519), .A3(net_3518), .A4(net_3517) );
SDFFS_X2 inst_2084 ( .QN(net_9057), .SI(net_6126), .SE(net_2946), .D(net_2912), .CK(net_11190), .SN(x6501) );
INV_X4 inst_5711 ( .A(net_8958), .ZN(net_1575) );
CLKBUF_X2 inst_16179 ( .A(net_16026), .Z(net_16027) );
CLKBUF_X2 inst_11534 ( .A(net_11381), .Z(net_11382) );
CLKBUF_X2 inst_12310 ( .A(net_12157), .Z(net_12158) );
CLKBUF_X2 inst_18715 ( .A(net_17559), .Z(net_18563) );
CLKBUF_X2 inst_17143 ( .A(net_16990), .Z(net_16991) );
AOI22_X2 inst_8203 ( .B1(net_8756), .A1(net_8386), .A2(net_3867), .B2(net_3866), .ZN(net_3833) );
CLKBUF_X2 inst_16686 ( .A(net_16533), .Z(net_16534) );
SDFF_X2 inst_803 ( .SI(net_8482), .Q(net_8482), .D(net_3961), .SE(net_3884), .CK(net_9985) );
CLKBUF_X2 inst_12011 ( .A(net_11858), .Z(net_11859) );
CLKBUF_X2 inst_18943 ( .A(net_18790), .Z(net_18791) );
CLKBUF_X2 inst_15167 ( .A(net_15014), .Z(net_15015) );
CLKBUF_X2 inst_10312 ( .A(net_9950), .Z(net_10160) );
CLKBUF_X2 inst_11936 ( .A(net_11783), .Z(net_11784) );
SDFF_X2 inst_662 ( .Q(net_8436), .D(net_8436), .SI(net_3953), .SE(net_3934), .CK(net_10252) );
CLKBUF_X2 inst_15590 ( .A(net_15273), .Z(net_15438) );
NOR2_X2 inst_3495 ( .A1(net_8217), .ZN(net_2222), .A2(net_2187) );
SDFF_X2 inst_1533 ( .Q(net_7881), .D(net_7881), .SI(net_2658), .SE(net_2543), .CK(net_15528) );
DFFR_X2 inst_7156 ( .QN(net_9054), .D(net_2854), .CK(net_11150), .RN(x6501) );
AOI22_X2 inst_7741 ( .B1(net_6970), .A1(net_6930), .ZN(net_5444), .A2(net_5443), .B2(net_5442) );
CLKBUF_X2 inst_11046 ( .A(net_9732), .Z(net_10894) );
CLKBUF_X2 inst_12491 ( .A(net_12338), .Z(net_12339) );
CLKBUF_X2 inst_17720 ( .A(net_17567), .Z(net_17568) );
CLKBUF_X2 inst_18574 ( .A(net_18421), .Z(net_18422) );
CLKBUF_X2 inst_18243 ( .A(net_18090), .Z(net_18091) );
CLKBUF_X2 inst_19050 ( .A(net_18897), .Z(net_18898) );
XOR2_X2 inst_53 ( .B(net_6839), .A(net_1029), .Z(net_994) );
INV_X8 inst_5030 ( .ZN(net_4364), .A(net_3351) );
CLKBUF_X2 inst_12653 ( .A(net_12500), .Z(net_12501) );
NOR2_X4 inst_3337 ( .ZN(net_2094), .A1(net_1890), .A2(net_1884) );
SDFFR_X2 inst_2614 ( .Q(net_7369), .D(net_7369), .SE(net_1136), .CK(net_18643), .RN(x6501), .SI(x4831) );
NAND2_X2 inst_4090 ( .ZN(net_5449), .A2(net_5252), .A1(net_5168) );
CLKBUF_X2 inst_10513 ( .A(net_9997), .Z(net_10361) );
SDFFR_X2 inst_2111 ( .SE(net_5582), .D(net_5525), .CK(net_14210), .RN(x6501), .SI(x76), .Q(x76) );
CLKBUF_X2 inst_14512 ( .A(net_14359), .Z(net_14360) );
AOI22_X2 inst_8419 ( .B1(net_6586), .A1(net_6553), .A2(net_6257), .B2(net_6110), .ZN(net_3523) );
CLKBUF_X2 inst_13943 ( .A(net_13790), .Z(net_13791) );
SDFF_X2 inst_1463 ( .SI(net_7287), .Q(net_7144), .D(net_7144), .SE(net_6279), .CK(net_14920) );
CLKBUF_X2 inst_14242 ( .A(net_14089), .Z(net_14090) );
CLKBUF_X2 inst_9665 ( .A(net_9512), .Z(net_9513) );
CLKBUF_X2 inst_16311 ( .A(net_15259), .Z(net_16159) );
CLKBUF_X2 inst_13463 ( .A(net_13310), .Z(net_13311) );
SDFF_X2 inst_759 ( .Q(net_8800), .D(net_8800), .SI(net_3963), .SE(net_3879), .CK(net_12334) );
CLKBUF_X2 inst_11655 ( .A(net_11153), .Z(net_11503) );
CLKBUF_X2 inst_13192 ( .A(net_11748), .Z(net_13040) );
CLKBUF_X2 inst_18776 ( .A(net_15815), .Z(net_18624) );
INV_X2 inst_6596 ( .A(net_6132), .ZN(net_6131) );
CLKBUF_X2 inst_9274 ( .A(net_9121), .Z(net_9122) );
CLKBUF_X2 inst_18330 ( .A(net_18177), .Z(net_18178) );
NOR2_X2 inst_3586 ( .ZN(net_1294), .A1(net_486), .A2(net_268) );
CLKBUF_X2 inst_13652 ( .A(net_13499), .Z(net_13500) );
AOI22_X2 inst_7744 ( .B1(net_6973), .A1(net_6933), .A2(net_5443), .B2(net_5442), .ZN(net_5430) );
CLKBUF_X2 inst_14625 ( .A(net_14472), .Z(net_14473) );
DFFR_X2 inst_7203 ( .D(net_2357), .QN(net_224), .CK(net_15008), .RN(x6501) );
CLKBUF_X2 inst_9974 ( .A(net_9821), .Z(net_9822) );
SDFFR_X2 inst_2282 ( .SE(net_2789), .SI(net_1330), .Q(net_254), .D(net_254), .CK(net_18331), .RN(x6501) );
CLKBUF_X2 inst_14594 ( .A(net_11638), .Z(net_14442) );
INV_X4 inst_5718 ( .A(net_8939), .ZN(net_2628) );
XNOR2_X2 inst_169 ( .ZN(net_1824), .A(net_1546), .B(net_1545) );
INV_X4 inst_6158 ( .ZN(net_6209), .A(net_6207) );
CLKBUF_X2 inst_12880 ( .A(net_12260), .Z(net_12728) );
CLKBUF_X2 inst_11748 ( .A(net_11595), .Z(net_11596) );
SDFF_X2 inst_555 ( .Q(net_8702), .D(net_8702), .SI(net_3949), .SE(net_3935), .CK(net_10564) );
AOI22_X2 inst_8014 ( .A1(net_7962), .B1(net_7792), .A2(net_6092), .B2(net_6091), .ZN(net_4121) );
CLKBUF_X2 inst_10293 ( .A(net_9204), .Z(net_10141) );
CLKBUF_X2 inst_12978 ( .A(net_9287), .Z(net_12826) );
SDFF_X2 inst_1184 ( .D(net_7316), .SI(net_6558), .Q(net_6558), .SE(net_3070), .CK(net_12066) );
CLKBUF_X2 inst_17148 ( .A(net_16995), .Z(net_16996) );
CLKBUF_X2 inst_9352 ( .A(net_9199), .Z(net_9200) );
NAND2_X2 inst_4685 ( .ZN(net_4385), .A1(net_2085), .A2(net_1913) );
CLKBUF_X2 inst_14325 ( .A(net_9325), .Z(net_14173) );
INV_X4 inst_6157 ( .A(net_6201), .ZN(net_6200) );
AOI22_X2 inst_7796 ( .B1(net_7183), .A2(net_6129), .B2(net_5655), .ZN(net_4793), .A1(net_1391) );
AOI22_X2 inst_8197 ( .B1(net_8792), .A1(net_8533), .A2(net_3861), .B2(net_3860), .ZN(net_3839) );
CLKBUF_X2 inst_12523 ( .A(net_12370), .Z(net_12371) );
CLKBUF_X2 inst_14999 ( .A(net_14277), .Z(net_14847) );
INV_X2 inst_6580 ( .A(net_5943), .ZN(x1152) );
CLKBUF_X2 inst_18754 ( .A(net_10723), .Z(net_18602) );
INV_X4 inst_5140 ( .ZN(net_3555), .A(net_3529) );
CLKBUF_X2 inst_9480 ( .A(net_9327), .Z(net_9328) );
CLKBUF_X2 inst_11863 ( .A(net_11710), .Z(net_11711) );
CLKBUF_X2 inst_11578 ( .A(net_9315), .Z(net_11426) );
AOI221_X2 inst_8756 ( .B2(net_5609), .ZN(net_5530), .A(net_5253), .C2(net_4388), .C1(net_2594), .B1(net_360) );
CLKBUF_X2 inst_12273 ( .A(net_12120), .Z(net_12121) );
DFFR_X1 inst_7521 ( .Q(net_7629), .D(net_1077), .CK(net_15714), .RN(x6501) );
AOI21_X2 inst_8952 ( .A(net_5783), .ZN(net_5664), .B1(net_5469), .B2(net_5263) );
CLKBUF_X2 inst_12931 ( .A(net_9753), .Z(net_12779) );
NAND3_X2 inst_3991 ( .A2(net_1925), .A3(net_1669), .ZN(net_1659), .A1(net_1591) );
CLKBUF_X2 inst_9546 ( .A(net_9393), .Z(net_9394) );
CLKBUF_X2 inst_13620 ( .A(net_13467), .Z(net_13468) );
CLKBUF_X2 inst_14812 ( .A(net_12379), .Z(net_14660) );
INV_X2 inst_6203 ( .ZN(net_5507), .A(net_5417) );
CLKBUF_X2 inst_15661 ( .A(net_13564), .Z(net_15509) );
NOR2_X2 inst_3343 ( .A2(net_6792), .ZN(net_5778), .A1(net_1912) );
AOI222_X1 inst_8617 ( .A2(net_8221), .ZN(net_4893), .A1(net_4891), .B2(net_4889), .C2(net_4888), .B1(net_4699), .C1(net_3108) );
NAND2_X2 inst_4140 ( .ZN(net_5380), .A1(net_5116), .A2(net_5115) );
CLKBUF_X2 inst_13340 ( .A(net_13187), .Z(net_13188) );
CLKBUF_X2 inst_16654 ( .A(net_16501), .Z(net_16502) );
OR3_X4 inst_2801 ( .A2(net_2965), .ZN(net_1434), .A1(net_1295), .A3(net_1294) );
NAND2_X2 inst_4219 ( .A1(net_6893), .A2(net_5247), .ZN(net_5241) );
SDFFR_X2 inst_2303 ( .D(net_7516), .SE(net_2748), .SI(net_432), .Q(net_432), .CK(net_13701), .RN(x6501) );
AND2_X2 inst_9153 ( .ZN(net_3090), .A2(net_3089), .A1(net_1066) );
CLKBUF_X2 inst_13714 ( .A(net_11267), .Z(net_13562) );
AOI22_X2 inst_8090 ( .B1(net_8176), .A1(net_7734), .B2(net_6101), .A2(net_6095), .ZN(net_4056) );
CLKBUF_X2 inst_14765 ( .A(net_14612), .Z(net_14613) );
CLKBUF_X2 inst_16991 ( .A(net_16838), .Z(net_16839) );
CLKBUF_X2 inst_16369 ( .A(net_16216), .Z(net_16217) );
NAND4_X2 inst_3771 ( .ZN(net_4250), .A1(net_3761), .A2(net_3760), .A3(net_3759), .A4(net_3758) );
CLKBUF_X2 inst_17895 ( .A(net_17742), .Z(net_17743) );
SDFF_X2 inst_1695 ( .SI(net_7856), .Q(net_7856), .D(net_2575), .SE(net_2558), .CK(net_15979) );
INV_X4 inst_5557 ( .ZN(net_631), .A(net_630) );
CLKBUF_X2 inst_17957 ( .A(net_17804), .Z(net_17805) );
AOI21_X2 inst_8954 ( .ZN(net_5592), .B2(net_5466), .B1(net_4923), .A(net_3386) );
CLKBUF_X2 inst_9724 ( .A(net_9571), .Z(net_9572) );
CLKBUF_X2 inst_15851 ( .A(net_15698), .Z(net_15699) );
SDFF_X2 inst_1339 ( .Q(net_7950), .D(net_7950), .SE(net_2755), .SI(net_2702), .CK(net_18873) );
NAND2_X2 inst_4284 ( .A1(net_7007), .A2(net_5249), .ZN(net_5176) );
CLKBUF_X2 inst_11235 ( .A(net_11082), .Z(net_11083) );
MUX2_X2 inst_4971 ( .A(net_6322), .Z(net_2068), .S(net_1700), .B(x4902) );
NAND2_X2 inst_4724 ( .A1(net_7374), .ZN(net_1974), .A2(net_1783) );
CLKBUF_X2 inst_17672 ( .A(net_13892), .Z(net_17520) );
NAND2_X2 inst_4467 ( .ZN(net_5022), .A2(net_4779), .A1(net_4508) );
CLKBUF_X2 inst_13512 ( .A(net_10197), .Z(net_13360) );
NAND4_X2 inst_3654 ( .A4(net_6036), .A1(net_6035), .ZN(net_4611), .A2(net_4168), .A3(net_4167) );
CLKBUF_X2 inst_18971 ( .A(net_18818), .Z(net_18819) );
SDFF_X2 inst_977 ( .SI(net_7313), .Q(net_6720), .D(net_6720), .SE(net_3124), .CK(net_12042) );
DFFS_X2 inst_6901 ( .Q(net_8214), .D(net_2257), .CK(net_17298), .SN(x6501) );
NAND2_X2 inst_4802 ( .ZN(net_5714), .A1(net_1136), .A2(net_575) );
XNOR2_X2 inst_297 ( .A(net_3138), .B(net_1468), .ZN(net_985) );
CLKBUF_X2 inst_15402 ( .A(net_15249), .Z(net_15250) );
CLKBUF_X2 inst_11728 ( .A(net_11575), .Z(net_11576) );
CLKBUF_X2 inst_13145 ( .A(net_12483), .Z(net_12993) );
CLKBUF_X2 inst_13933 ( .A(net_13780), .Z(net_13781) );
CLKBUF_X2 inst_16334 ( .A(net_16181), .Z(net_16182) );
NOR2_X2 inst_3436 ( .A1(net_7650), .A2(net_3081), .ZN(net_3073) );
SDFFR_X2 inst_2188 ( .QN(net_7218), .SI(net_2981), .D(net_2798), .SE(net_1379), .CK(net_15149), .RN(x6501) );
NOR2_X2 inst_3351 ( .ZN(net_5574), .A1(net_5424), .A2(net_5423) );
CLKBUF_X2 inst_10466 ( .A(net_10313), .Z(net_10314) );
CLKBUF_X2 inst_13057 ( .A(net_12904), .Z(net_12905) );
CLKBUF_X2 inst_17692 ( .A(net_17539), .Z(net_17540) );
XNOR2_X2 inst_162 ( .B(net_7653), .ZN(net_1845), .A(net_1569) );
CLKBUF_X2 inst_17645 ( .A(net_17492), .Z(net_17493) );
NOR3_X2 inst_3308 ( .ZN(net_1566), .A1(net_1565), .A2(net_530), .A3(x13884) );
DFFR_X1 inst_7373 ( .QN(net_5945), .D(net_5888), .CK(net_9408), .RN(x6501) );
CLKBUF_X2 inst_14903 ( .A(net_14750), .Z(net_14751) );
DFFR_X2 inst_7302 ( .D(net_6479), .QN(net_6476), .CK(net_11729), .RN(x6501) );
CLKBUF_X2 inst_17697 ( .A(net_17544), .Z(net_17545) );
CLKBUF_X2 inst_13387 ( .A(net_13234), .Z(net_13235) );
NAND4_X2 inst_3819 ( .ZN(net_3607), .A1(net_3411), .A2(net_3410), .A3(net_3409), .A4(net_3408) );
OR2_X4 inst_2829 ( .ZN(net_3529), .A1(net_3359), .A2(net_3301) );
CLKBUF_X2 inst_15939 ( .A(net_15786), .Z(net_15787) );
CLKBUF_X2 inst_18902 ( .A(net_18574), .Z(net_18750) );
NAND4_X2 inst_3668 ( .A4(net_6044), .A1(net_6043), .ZN(net_4597), .A2(net_4084), .A3(net_4083) );
CLKBUF_X2 inst_11383 ( .A(net_11230), .Z(net_11231) );
CLKBUF_X2 inst_16790 ( .A(net_15958), .Z(net_16638) );
CLKBUF_X2 inst_12086 ( .A(net_11933), .Z(net_11934) );
AOI22_X2 inst_8143 ( .B1(net_8119), .A1(net_7881), .A2(net_6098), .B2(net_4190), .ZN(net_4008) );
CLKBUF_X2 inst_17681 ( .A(net_17528), .Z(net_17529) );
SDFF_X2 inst_1098 ( .D(net_7326), .SI(net_6535), .Q(net_6535), .SE(net_3086), .CK(net_11281) );
NAND2_X2 inst_4149 ( .ZN(net_5368), .A1(net_5107), .A2(net_5106) );
DFFR_X2 inst_7077 ( .Q(net_6346), .D(net_3876), .CK(net_17637), .RN(x6501) );
SDFFR_X2 inst_2443 ( .SE(net_2685), .D(net_2668), .SI(net_445), .Q(net_445), .CK(net_13827), .RN(x6501) );
CLKBUF_X2 inst_10051 ( .A(net_9898), .Z(net_9899) );
SDFF_X2 inst_723 ( .SI(net_8486), .Q(net_8486), .D(net_3938), .SE(net_3884), .CK(net_13032) );
AOI21_X2 inst_8921 ( .B2(net_5871), .ZN(net_5709), .A(net_5700), .B1(net_2728) );
CLKBUF_X2 inst_10990 ( .A(net_10837), .Z(net_10838) );
NAND3_X2 inst_3893 ( .ZN(net_5645), .A1(net_5574), .A3(net_5508), .A2(net_5422) );
CLKBUF_X2 inst_11055 ( .A(net_10698), .Z(net_10903) );
CLKBUF_X2 inst_11616 ( .A(net_11463), .Z(net_11464) );
INV_X4 inst_5777 ( .A(net_7564), .ZN(net_554) );
CLKBUF_X2 inst_13274 ( .A(net_12183), .Z(net_13122) );
CLKBUF_X2 inst_18836 ( .A(net_18683), .Z(net_18684) );
SDFFS_X2 inst_2067 ( .SI(net_2796), .SE(net_2417), .Q(net_180), .D(net_180), .CK(net_14943), .SN(x6501) );
AOI22_X2 inst_7894 ( .B1(net_8975), .A2(net_5538), .B2(net_5456), .ZN(net_4535), .A1(net_404) );
CLKBUF_X2 inst_14651 ( .A(net_14498), .Z(net_14499) );
CLKBUF_X2 inst_18018 ( .A(net_17865), .Z(net_17866) );
CLKBUF_X2 inst_17851 ( .A(net_17029), .Z(net_17699) );
AOI22_X2 inst_8268 ( .B1(net_8690), .A1(net_8653), .B2(net_6109), .A2(net_3857), .ZN(net_3770) );
CLKBUF_X2 inst_13075 ( .A(net_12922), .Z(net_12923) );
SDFFR_X1 inst_2777 ( .D(net_7388), .Q(net_7285), .SI(net_1946), .SE(net_1327), .CK(net_18168), .RN(x6501) );
CLKBUF_X2 inst_12283 ( .A(net_12130), .Z(net_12131) );
DFF_X1 inst_6784 ( .Q(net_7533), .D(net_4586), .CK(net_9390) );
DFF_X1 inst_6830 ( .Q(net_6450), .D(net_3618), .CK(net_15172) );
CLKBUF_X2 inst_17031 ( .A(net_16878), .Z(net_16879) );
CLKBUF_X2 inst_18360 ( .A(net_18207), .Z(net_18208) );
SDFFR_X2 inst_2446 ( .D(net_3056), .SE(net_2313), .SI(net_412), .Q(net_412), .CK(net_13933), .RN(x6501) );
INV_X8 inst_5046 ( .A(net_6126), .ZN(net_6124) );
CLKBUF_X2 inst_13602 ( .A(net_13449), .Z(net_13450) );
AOI22_X2 inst_7840 ( .A2(net_5595), .ZN(net_4670), .B1(net_4669), .B2(net_4388), .A1(net_310) );
AOI22_X2 inst_8452 ( .B1(net_6537), .A1(net_6504), .A2(net_6137), .B2(net_6104), .ZN(net_3488) );
CLKBUF_X2 inst_19094 ( .A(net_18941), .Z(net_18942) );
CLKBUF_X2 inst_14128 ( .A(net_10257), .Z(net_13976) );
CLKBUF_X2 inst_13070 ( .A(net_9905), .Z(net_12918) );
CLKBUF_X2 inst_15549 ( .A(net_15396), .Z(net_15397) );
CLKBUF_X2 inst_14260 ( .A(net_10862), .Z(net_14108) );
INV_X4 inst_5210 ( .ZN(net_2683), .A(net_2220) );
INV_X2 inst_6613 ( .A(net_7415), .ZN(net_6204) );
CLKBUF_X2 inst_12767 ( .A(net_12614), .Z(net_12615) );
CLKBUF_X2 inst_17820 ( .A(net_17667), .Z(net_17668) );
CLKBUF_X2 inst_16611 ( .A(net_12213), .Z(net_16459) );
INV_X4 inst_5464 ( .A(net_1810), .ZN(net_761) );
CLKBUF_X2 inst_16676 ( .A(net_16523), .Z(net_16524) );
CLKBUF_X2 inst_18718 ( .A(net_10135), .Z(net_18566) );
CLKBUF_X2 inst_14089 ( .A(net_12583), .Z(net_13937) );
CLKBUF_X2 inst_18070 ( .A(net_12299), .Z(net_17918) );
CLKBUF_X2 inst_18438 ( .A(net_18285), .Z(net_18286) );
AOI22_X2 inst_8366 ( .B1(net_8703), .A1(net_8666), .B2(net_6109), .A2(net_3857), .ZN(net_3682) );
SDFF_X2 inst_1818 ( .D(net_7275), .SI(net_7012), .Q(net_7012), .SE(net_6277), .CK(net_17367) );
DFFR_X2 inst_7110 ( .QN(net_7309), .D(net_3150), .CK(net_9654), .RN(x6501) );
CLKBUF_X2 inst_18341 ( .A(net_14676), .Z(net_18189) );
CLKBUF_X2 inst_10705 ( .A(net_10552), .Z(net_10553) );
CLKBUF_X2 inst_14706 ( .A(net_14553), .Z(net_14554) );
CLKBUF_X2 inst_10264 ( .A(net_10111), .Z(net_10112) );
SDFF_X2 inst_1766 ( .D(net_7283), .SI(net_6860), .Q(net_6860), .SE(net_6282), .CK(net_19020) );
CLKBUF_X2 inst_13888 ( .A(net_13735), .Z(net_13736) );
CLKBUF_X2 inst_18897 ( .A(net_9753), .Z(net_18745) );
AOI22_X2 inst_8216 ( .B1(net_8832), .A1(net_8351), .A2(net_6265), .B2(net_6253), .ZN(net_3820) );
CLKBUF_X2 inst_15398 ( .A(net_15245), .Z(net_15246) );
CLKBUF_X2 inst_9639 ( .A(net_9179), .Z(net_9487) );
NAND2_X2 inst_4548 ( .A1(net_3373), .ZN(net_3316), .A2(net_3315) );
CLKBUF_X2 inst_17679 ( .A(net_15638), .Z(net_17527) );
SDFF_X2 inst_876 ( .Q(net_8587), .D(net_8587), .SI(net_3951), .SE(net_3878), .CK(net_10593) );
OAI21_X4 inst_2979 ( .ZN(net_6145), .B1(net_4926), .A(net_3324), .B2(net_2161) );
NAND2_X2 inst_4727 ( .A1(net_7366), .ZN(net_2054), .A2(net_1782) );
CLKBUF_X2 inst_19182 ( .A(net_19029), .Z(net_19030) );
SDFFR_X2 inst_2433 ( .D(net_3334), .SE(net_2313), .SI(net_424), .Q(net_424), .CK(net_14547), .RN(x6501) );
CLKBUF_X2 inst_11665 ( .A(net_11512), .Z(net_11513) );
CLKBUF_X2 inst_11751 ( .A(net_11598), .Z(net_11599) );
SDFFR_X2 inst_2480 ( .Q(net_8990), .D(net_8990), .SI(net_4522), .SE(net_2562), .CK(net_13923), .RN(x6501) );
SDFF_X2 inst_562 ( .Q(net_8815), .D(net_8815), .SE(net_3964), .SI(net_3961), .CK(net_10165) );
CLKBUF_X2 inst_9845 ( .A(net_9572), .Z(net_9693) );
AOI21_X2 inst_8917 ( .ZN(net_5758), .A(net_5745), .B2(net_5594), .B1(net_4790) );
CLKBUF_X2 inst_14714 ( .A(net_13989), .Z(net_14562) );
INV_X2 inst_6385 ( .ZN(net_1321), .A(net_1320) );
CLKBUF_X2 inst_11445 ( .A(net_11292), .Z(net_11293) );
CLKBUF_X2 inst_15006 ( .A(net_14853), .Z(net_14854) );
AOI22_X2 inst_8277 ( .B1(net_8840), .A1(net_8359), .A2(net_6265), .B2(net_6253), .ZN(net_3764) );
MUX2_X2 inst_4953 ( .A(net_7385), .Z(net_2371), .S(net_2370), .B(net_798) );
CLKBUF_X2 inst_12404 ( .A(net_12251), .Z(net_12252) );
CLKBUF_X2 inst_9589 ( .A(net_9110), .Z(net_9437) );
DFFR_X2 inst_7164 ( .QN(net_8946), .D(net_2654), .CK(net_16314), .RN(x6501) );
NAND4_X2 inst_3659 ( .A4(net_6010), .A1(net_6009), .ZN(net_4606), .A2(net_4138), .A3(net_4137) );
NOR2_X2 inst_3604 ( .ZN(net_2762), .A1(net_1057), .A2(net_833) );
DFFR_X1 inst_7465 ( .QN(net_7433), .D(net_4378), .CK(net_10121), .RN(x6501) );
CLKBUF_X2 inst_17028 ( .A(net_16875), .Z(net_16876) );
SDFF_X2 inst_1109 ( .D(net_7313), .SI(net_6522), .Q(net_6522), .SE(net_3086), .CK(net_12001) );
INV_X2 inst_6487 ( .A(net_6350), .ZN(net_2079) );
CLKBUF_X2 inst_12054 ( .A(net_9587), .Z(net_11902) );
OAI21_X2 inst_3037 ( .B2(net_8237), .B1(net_4928), .ZN(net_4841), .A(net_3237) );
CLKBUF_X2 inst_11522 ( .A(net_11369), .Z(net_11370) );
CLKBUF_X2 inst_14857 ( .A(net_14704), .Z(net_14705) );
SDFF_X2 inst_1314 ( .SI(net_7675), .Q(net_7675), .SE(net_2714), .D(net_2659), .CK(net_15540) );
AOI22_X2 inst_7956 ( .B1(net_8091), .A1(net_7751), .B2(net_6108), .A2(net_6096), .ZN(net_4171) );
SDFF_X2 inst_1156 ( .SI(net_7339), .Q(net_6614), .D(net_6614), .SE(net_3069), .CK(net_11861) );
INV_X4 inst_5533 ( .A(net_669), .ZN(net_656) );
NOR2_X2 inst_3378 ( .ZN(net_5547), .A1(net_5313), .A2(net_5312) );
CLKBUF_X2 inst_11466 ( .A(net_11313), .Z(net_11314) );
CLKBUF_X2 inst_16458 ( .A(net_16305), .Z(net_16306) );
INV_X4 inst_5993 ( .A(net_6292), .ZN(net_2673) );
CLKBUF_X2 inst_12512 ( .A(net_12359), .Z(net_12360) );
CLKBUF_X2 inst_13676 ( .A(net_13523), .Z(net_13524) );
CLKBUF_X2 inst_14259 ( .A(net_12796), .Z(net_14107) );
SDFF_X2 inst_1880 ( .D(net_7290), .SI(net_6987), .Q(net_6987), .SE(net_6283), .CK(net_15322) );
SDFF_X2 inst_1295 ( .Q(net_8099), .D(net_8099), .SI(net_2713), .SE(net_2707), .CK(net_13789) );
DFFR_X1 inst_7457 ( .Q(net_7163), .D(net_4727), .CK(net_9599), .RN(x6501) );
XNOR2_X2 inst_262 ( .B(net_8894), .ZN(net_1168), .A(net_1167) );
NAND4_X2 inst_3630 ( .ZN(net_5540), .A2(net_5280), .A1(net_5047), .A3(net_4659), .A4(net_4570) );
NAND2_X2 inst_4675 ( .A2(net_7485), .ZN(net_2296), .A1(net_2112) );
CLKBUF_X2 inst_10333 ( .A(net_10180), .Z(net_10181) );
CLKBUF_X2 inst_16644 ( .A(net_16491), .Z(net_16492) );
SDFF_X2 inst_1035 ( .SI(net_7342), .Q(net_6716), .D(net_6716), .SE(net_3125), .CK(net_11682) );
AOI22_X2 inst_7942 ( .B1(net_7919), .A1(net_7817), .B2(net_6103), .A2(net_4398), .ZN(net_4183) );
CLKBUF_X2 inst_18466 ( .A(net_12598), .Z(net_18314) );
NAND4_X2 inst_3637 ( .ZN(net_5253), .A4(net_4793), .A1(net_4693), .A3(net_4692), .A2(net_4572) );
CLKBUF_X2 inst_11490 ( .A(net_11337), .Z(net_11338) );
CLKBUF_X2 inst_17286 ( .A(net_17133), .Z(net_17134) );
SDFF_X2 inst_1883 ( .D(net_7294), .SI(net_6991), .Q(net_6991), .SE(net_6283), .CK(net_17668) );
DFFR_X2 inst_7240 ( .QN(net_6751), .D(net_2209), .CK(net_17930), .RN(x6501) );
CLKBUF_X2 inst_9580 ( .A(net_9427), .Z(net_9428) );
CLKBUF_X2 inst_12863 ( .A(net_12710), .Z(net_12711) );
NOR2_X1 inst_3621 ( .A2(net_4371), .ZN(net_2000), .A1(net_1656) );
SDFF_X2 inst_864 ( .Q(net_8573), .D(net_8573), .SI(net_3967), .SE(net_3878), .CK(net_12241) );
XOR2_X1 inst_86 ( .Z(net_2034), .B(net_2033), .A(net_1767) );
SDFF_X2 inst_949 ( .SI(net_7332), .Q(net_6706), .D(net_6706), .SE(net_3125), .CK(net_9085) );
CLKBUF_X2 inst_18306 ( .A(net_11206), .Z(net_18154) );
NOR3_X2 inst_3283 ( .A1(net_2400), .ZN(net_2320), .A3(net_2317), .A2(net_1770) );
CLKBUF_X2 inst_12580 ( .A(net_12427), .Z(net_12428) );
CLKBUF_X2 inst_16195 ( .A(net_16042), .Z(net_16043) );
CLKBUF_X2 inst_15651 ( .A(net_15498), .Z(net_15499) );
NAND4_X2 inst_3730 ( .ZN(net_4300), .A1(net_4136), .A2(net_4135), .A3(net_4134), .A4(net_4133) );
CLKBUF_X2 inst_13294 ( .A(net_12138), .Z(net_13142) );
NOR2_X2 inst_3598 ( .ZN(net_1162), .A1(net_1011), .A2(net_845) );
CLKBUF_X2 inst_10342 ( .A(net_10189), .Z(net_10190) );
CLKBUF_X2 inst_17237 ( .A(net_17084), .Z(net_17085) );
SDFFR_X2 inst_2109 ( .SI(net_7409), .Q(net_7409), .SE(net_6198), .D(net_5731), .CK(net_9377), .RN(x6501) );
SDFF_X2 inst_1826 ( .D(net_7279), .SI(net_6856), .Q(net_6856), .SE(net_6282), .CK(net_14626) );
CLKBUF_X2 inst_12140 ( .A(net_10920), .Z(net_11988) );
INV_X4 inst_5395 ( .A(net_1138), .ZN(net_1049) );
SDFF_X2 inst_2020 ( .SI(net_7922), .Q(net_7922), .D(net_2589), .SE(net_2461), .CK(net_15564) );
INV_X2 inst_6192 ( .A(net_6787), .ZN(net_5734) );
NAND2_X2 inst_4361 ( .A1(net_7070), .A2(net_5162), .ZN(net_5096) );
OR2_X4 inst_2820 ( .A1(net_6164), .ZN(net_4954), .A2(net_4387) );
CLKBUF_X2 inst_13721 ( .A(net_13568), .Z(net_13569) );
SDFFR_X2 inst_2404 ( .D(net_7368), .SE(net_2734), .SI(net_274), .Q(net_274), .CK(net_13680), .RN(x6501) );
CLKBUF_X2 inst_14417 ( .A(net_14264), .Z(net_14265) );
AOI22_X2 inst_7994 ( .B1(net_8165), .A1(net_7723), .B2(net_6101), .A2(net_6095), .ZN(net_6010) );
CLKBUF_X2 inst_14075 ( .A(net_13922), .Z(net_13923) );
CLKBUF_X2 inst_15539 ( .A(net_15386), .Z(net_15387) );
SDFF_X2 inst_1578 ( .Q(net_8011), .D(net_8011), .SI(net_2585), .SE(net_2545), .CK(net_18550) );
AOI22_X2 inst_7849 ( .A2(net_5595), .ZN(net_4659), .B2(net_4388), .B1(net_2616), .A1(net_318) );
CLKBUF_X2 inst_17714 ( .A(net_17561), .Z(net_17562) );
AND2_X4 inst_9053 ( .ZN(net_3573), .A1(net_3359), .A2(net_3358) );
NAND2_X2 inst_4612 ( .A2(net_6144), .ZN(net_2617), .A1(net_2616) );
CLKBUF_X2 inst_9598 ( .A(net_9445), .Z(net_9446) );
CLKBUF_X2 inst_11398 ( .A(net_11245), .Z(net_11246) );
CLKBUF_X2 inst_15676 ( .A(net_15523), .Z(net_15524) );
AOI221_X2 inst_8820 ( .C1(net_7181), .B2(net_6432), .C2(net_5655), .B1(net_5654), .A(net_4905), .ZN(net_4678) );
CLKBUF_X2 inst_18802 ( .A(net_18649), .Z(net_18650) );
XNOR2_X2 inst_175 ( .B(net_2669), .ZN(net_1765), .A(net_1677) );
CLKBUF_X2 inst_11989 ( .A(net_9154), .Z(net_11837) );
INV_X8 inst_5010 ( .ZN(net_4708), .A(net_4455) );
CLKBUF_X2 inst_10491 ( .A(net_10338), .Z(net_10339) );
CLKBUF_X2 inst_18596 ( .A(net_18443), .Z(net_18444) );
CLKBUF_X2 inst_15764 ( .A(net_15611), .Z(net_15612) );
SDFF_X2 inst_1737 ( .SI(net_7297), .Q(net_7154), .D(net_7154), .SE(net_6279), .CK(net_18191) );
CLKBUF_X2 inst_10895 ( .A(net_10742), .Z(net_10743) );
OAI21_X2 inst_2995 ( .B2(net_5902), .ZN(net_5898), .A(net_5829), .B1(net_614) );
AOI222_X1 inst_8594 ( .B2(net_6763), .ZN(net_5851), .B1(net_5835), .A2(net_5832), .C2(net_5824), .C1(net_2121), .A1(x3327) );
DFFR_X2 inst_7081 ( .QN(net_7665), .D(net_3892), .CK(net_12684), .RN(x6501) );
INV_X4 inst_5513 ( .ZN(net_3241), .A(net_680) );
NAND2_X2 inst_4541 ( .A1(net_3374), .A2(net_3369), .ZN(net_3365) );
CLKBUF_X2 inst_14073 ( .A(net_13920), .Z(net_13921) );
CLKBUF_X2 inst_18017 ( .A(net_16243), .Z(net_17865) );
SDFF_X2 inst_1149 ( .SI(net_7330), .Q(net_6605), .D(net_6605), .SE(net_3069), .CK(net_11278) );
CLKBUF_X2 inst_10146 ( .A(net_9370), .Z(net_9994) );
CLKBUF_X2 inst_14354 ( .A(net_14201), .Z(net_14202) );
INV_X4 inst_5640 ( .A(net_7432), .ZN(net_3581) );
CLKBUF_X2 inst_9696 ( .A(net_9176), .Z(net_9544) );
CLKBUF_X2 inst_11475 ( .A(net_9990), .Z(net_11323) );
NAND2_X2 inst_4719 ( .A1(net_7370), .ZN(net_1977), .A2(net_1784) );
CLKBUF_X2 inst_15026 ( .A(net_14873), .Z(net_14874) );
CLKBUF_X2 inst_17617 ( .A(net_15280), .Z(net_17465) );
NAND2_X2 inst_4353 ( .A1(net_7149), .A2(net_5166), .ZN(net_5104) );
INV_X4 inst_6003 ( .ZN(net_2634), .A(net_158) );
CLKBUF_X2 inst_9285 ( .A(net_9132), .Z(net_9133) );
NAND3_X2 inst_3934 ( .ZN(net_5516), .A1(net_5278), .A2(net_4656), .A3(net_4567) );
CLKBUF_X2 inst_9716 ( .A(net_9328), .Z(net_9564) );
CLKBUF_X2 inst_17602 ( .A(net_17449), .Z(net_17450) );
SDFF_X2 inst_948 ( .SI(net_7312), .Q(net_6686), .D(net_6686), .SE(net_3125), .CK(net_12052) );
CLKBUF_X2 inst_12475 ( .A(net_11229), .Z(net_12323) );
CLKBUF_X2 inst_13302 ( .A(net_13149), .Z(net_13150) );
CLKBUF_X2 inst_17250 ( .A(net_17097), .Z(net_17098) );
CLKBUF_X2 inst_18414 ( .A(net_18261), .Z(net_18262) );
CLKBUF_X2 inst_14795 ( .A(net_14642), .Z(net_14643) );
INV_X16 inst_6644 ( .ZN(net_3879), .A(net_3307) );
CLKBUF_X2 inst_13493 ( .A(net_13340), .Z(net_13341) );
CLKBUF_X2 inst_11407 ( .A(net_11254), .Z(net_11255) );
CLKBUF_X2 inst_16079 ( .A(net_12353), .Z(net_15927) );
CLKBUF_X2 inst_11275 ( .A(net_11122), .Z(net_11123) );
CLKBUF_X2 inst_15892 ( .A(net_9982), .Z(net_15740) );
AOI22_X2 inst_8039 ( .B1(net_8136), .A1(net_7898), .A2(net_6098), .B2(net_4190), .ZN(net_4100) );
CLKBUF_X2 inst_11647 ( .A(net_10799), .Z(net_11495) );
CLKBUF_X2 inst_15579 ( .A(net_15426), .Z(net_15427) );
INV_X4 inst_5444 ( .ZN(net_2571), .A(net_816) );
CLKBUF_X2 inst_9966 ( .A(net_9813), .Z(net_9814) );
CLKBUF_X2 inst_14671 ( .A(net_14518), .Z(net_14519) );
SDFF_X2 inst_2002 ( .SI(net_7791), .Q(net_7791), .D(net_2722), .SE(net_2459), .CK(net_15950) );
NAND2_X2 inst_4380 ( .A1(net_7157), .A2(net_5166), .ZN(net_5077) );
INV_X4 inst_6030 ( .A(net_6376), .ZN(net_504) );
AOI22_X2 inst_8430 ( .B1(net_6664), .A1(net_6631), .A2(net_6213), .B2(net_6138), .ZN(net_3511) );
CLKBUF_X2 inst_10471 ( .A(net_10318), .Z(net_10319) );
SDFF_X2 inst_608 ( .SI(net_8403), .Q(net_8403), .SE(net_3969), .D(net_3950), .CK(net_10548) );
SDFF_X2 inst_834 ( .SI(net_8643), .Q(net_8643), .D(net_3966), .SE(net_3885), .CK(net_10893) );
CLKBUF_X2 inst_11183 ( .A(net_10052), .Z(net_11031) );
CLKBUF_X2 inst_16869 ( .A(net_16716), .Z(net_16717) );
OAI22_X2 inst_2920 ( .ZN(net_3191), .B1(net_3190), .A2(net_3163), .B2(net_2767), .A1(net_1140) );
AOI221_X4 inst_8729 ( .B1(net_8706), .C1(net_8484), .B2(net_4350), .C2(net_4349), .ZN(net_4336), .A(net_4245) );
SDFF_X2 inst_966 ( .SI(net_7326), .Q(net_6733), .D(net_6733), .SE(net_3124), .CK(net_11300) );
CLKBUF_X2 inst_14951 ( .A(net_10548), .Z(net_14799) );
OAI221_X2 inst_2961 ( .B1(net_7173), .ZN(net_4553), .C2(net_4401), .C1(net_4385), .A(net_4320), .B2(net_2106) );
DFFR_X2 inst_7189 ( .QN(net_6317), .D(net_2470), .CK(net_14823), .RN(x6501) );
AOI21_X2 inst_8924 ( .B2(net_5871), .ZN(net_5699), .A(net_5698), .B1(x552) );
CLKBUF_X2 inst_11833 ( .A(net_10961), .Z(net_11681) );
SDFFR_X2 inst_2506 ( .Q(net_8999), .D(net_8999), .SI(net_2600), .SE(net_2562), .CK(net_14695), .RN(x6501) );
CLKBUF_X2 inst_13214 ( .A(net_13061), .Z(net_13062) );
INV_X4 inst_5836 ( .A(net_7259), .ZN(net_1994) );
INV_X4 inst_5976 ( .A(net_7443), .ZN(net_3921) );
INV_X4 inst_5245 ( .ZN(net_5582), .A(net_1822) );
INV_X4 inst_5575 ( .A(net_6324), .ZN(net_1639) );
NAND2_X2 inst_4557 ( .A1(net_6386), .A2(net_6184), .ZN(net_3253) );
NOR2_X2 inst_3607 ( .ZN(net_1067), .A2(net_845), .A1(net_555) );
AOI22_X2 inst_8583 ( .B2(net_6318), .ZN(net_1794), .B1(net_1254), .A2(net_636), .A1(x4392) );
CLKBUF_X2 inst_10498 ( .A(net_10345), .Z(net_10346) );
CLKBUF_X2 inst_13324 ( .A(net_13171), .Z(net_13172) );
CLKBUF_X2 inst_16395 ( .A(net_11620), .Z(net_16243) );
OAI21_X2 inst_3160 ( .B2(net_2304), .ZN(net_1926), .B1(net_1925), .A(net_1591) );
CLKBUF_X2 inst_14022 ( .A(net_11762), .Z(net_13870) );
OR2_X4 inst_2861 ( .ZN(net_6282), .A1(net_2200), .A2(net_2199) );
CLKBUF_X2 inst_14825 ( .A(net_14672), .Z(net_14673) );
XOR2_X2 inst_66 ( .A(net_6320), .B(net_6319), .Z(net_797) );
NAND2_X2 inst_4814 ( .A2(net_2520), .ZN(net_1255), .A1(x3762) );
CLKBUF_X2 inst_11139 ( .A(net_10772), .Z(net_10987) );
CLKBUF_X2 inst_11012 ( .A(net_10859), .Z(net_10860) );
AOI22_X2 inst_7920 ( .A1(net_8982), .A2(net_5456), .B2(net_5260), .ZN(net_4462), .B1(net_2916) );
CLKBUF_X2 inst_10604 ( .A(net_10451), .Z(net_10452) );
AOI221_X2 inst_8807 ( .C2(net_5535), .A(net_5520), .B2(net_5260), .ZN(net_4721), .B1(net_3388), .C1(net_469) );
XNOR2_X2 inst_273 ( .A(net_2936), .ZN(net_1040), .B(net_1039) );
CLKBUF_X2 inst_12297 ( .A(net_12144), .Z(net_12145) );
CLKBUF_X2 inst_13443 ( .A(net_12703), .Z(net_13291) );
CLKBUF_X2 inst_15365 ( .A(net_15212), .Z(net_15213) );
SDFFR_X2 inst_2418 ( .D(net_2686), .SE(net_2685), .SI(net_464), .Q(net_464), .CK(net_16914), .RN(x6501) );
SDFF_X2 inst_366 ( .SI(net_8331), .Q(net_8331), .SE(net_3978), .D(net_3939), .CK(net_12568) );
INV_X4 inst_6162 ( .A(net_6272), .ZN(net_6267) );
DFFR_X2 inst_7019 ( .QN(net_6301), .D(net_5692), .CK(net_16939), .RN(x6501) );
CLKBUF_X2 inst_9397 ( .A(net_9244), .Z(net_9245) );
CLKBUF_X2 inst_9565 ( .A(net_9244), .Z(net_9413) );
CLKBUF_X2 inst_12542 ( .A(net_12389), .Z(net_12390) );
AOI22_X2 inst_7964 ( .B1(net_8160), .A1(net_7718), .B2(net_6101), .A2(net_6095), .ZN(net_4164) );
CLKBUF_X2 inst_16845 ( .A(net_12091), .Z(net_16693) );
CLKBUF_X2 inst_16737 ( .A(net_16584), .Z(net_16585) );
DFFR_X2 inst_7313 ( .D(net_295), .QN(net_154), .CK(net_11133), .RN(x6501) );
NAND2_X2 inst_4746 ( .ZN(net_2574), .A2(net_1586), .A1(net_1023) );
INV_X4 inst_5896 ( .ZN(net_1058), .A(x12843) );
AOI22_X2 inst_7950 ( .B1(net_8022), .A1(net_7988), .B2(net_6102), .A2(net_6097), .ZN(net_4176) );
CLKBUF_X2 inst_18353 ( .A(net_11644), .Z(net_18201) );
SDFF_X2 inst_707 ( .SI(net_8624), .Q(net_8624), .SE(net_3984), .D(net_3951), .CK(net_13402) );
SDFF_X2 inst_1025 ( .SI(net_7332), .Q(net_6739), .D(net_6739), .SE(net_3124), .CK(net_9429) );
NAND2_X2 inst_4655 ( .A1(net_2700), .A2(net_2334), .ZN(net_2273) );
NAND4_X2 inst_3670 ( .A4(net_6046), .A1(net_6045), .ZN(net_4595), .A2(net_4072), .A3(net_4071) );
DFFR_X1 inst_7566 ( .Q(net_6826), .D(net_6814), .CK(net_18664), .RN(x6501) );
DFFR_X1 inst_7570 ( .D(net_6406), .QN(net_6405), .CK(net_9659), .RN(x6501) );
INV_X4 inst_5635 ( .A(net_7388), .ZN(net_922) );
AOI22_X2 inst_7834 ( .A2(net_6428), .B2(net_5657), .A1(net_5654), .ZN(net_4687), .B1(net_2731) );
INV_X4 inst_5542 ( .ZN(net_646), .A(x3762) );
AOI222_X1 inst_8654 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3912), .C1(net_1444), .B1(net_1314), .A1(x13921) );
CLKBUF_X2 inst_10080 ( .A(net_9927), .Z(net_9928) );
CLKBUF_X2 inst_16730 ( .A(net_10333), .Z(net_16578) );
CLKBUF_X2 inst_15094 ( .A(net_14941), .Z(net_14942) );
SDFFR_X2 inst_2576 ( .D(net_7393), .QN(net_7253), .SI(net_1960), .SE(net_1379), .CK(net_18321), .RN(x6501) );
DFFR_X2 inst_7269 ( .QN(net_7233), .D(net_1989), .CK(net_14778), .RN(x6501) );
CLKBUF_X2 inst_13654 ( .A(net_13501), .Z(net_13502) );
CLKBUF_X2 inst_13710 ( .A(net_13557), .Z(net_13558) );
SDFFR_X2 inst_2631 ( .Q(net_7392), .D(net_7392), .SE(net_1136), .CK(net_15795), .RN(x6501), .SI(x4503) );
CLKBUF_X2 inst_15988 ( .A(net_15835), .Z(net_15836) );
NAND4_X2 inst_3810 ( .ZN(net_3616), .A1(net_3447), .A2(net_3446), .A3(net_3445), .A4(net_3444) );
AOI22_X2 inst_8453 ( .B1(net_6736), .A1(net_6703), .B2(net_6202), .A2(net_3520), .ZN(net_3487) );
CLKBUF_X2 inst_13261 ( .A(net_11006), .Z(net_13109) );
NAND2_X2 inst_4523 ( .A2(net_3568), .ZN(net_3567), .A1(net_3566) );
DFFR_X2 inst_7073 ( .QN(net_8898), .D(net_4227), .CK(net_13530), .RN(x6501) );
SDFFR_X2 inst_2636 ( .Q(net_7375), .D(net_7375), .SE(net_1136), .CK(net_18604), .RN(x6501), .SI(x4778) );
INV_X2 inst_6198 ( .ZN(net_5512), .A(net_5437) );
CLKBUF_X2 inst_18039 ( .A(net_17886), .Z(net_17887) );
DFFR_X2 inst_7186 ( .QN(net_8961), .D(net_2492), .CK(net_15069), .RN(x6501) );
CLKBUF_X2 inst_16380 ( .A(net_16227), .Z(net_16228) );
DFFR_X1 inst_7579 ( .Q(net_393), .D(net_268), .CK(net_10808), .RN(x6501) );
CLKBUF_X2 inst_16038 ( .A(net_15265), .Z(net_15886) );
CLKBUF_X2 inst_11561 ( .A(net_10035), .Z(net_11409) );
CLKBUF_X2 inst_14491 ( .A(net_14338), .Z(net_14339) );
SDFF_X2 inst_445 ( .Q(net_8775), .D(net_8775), .SE(net_3982), .SI(net_3939), .CK(net_10580) );
CLKBUF_X2 inst_12961 ( .A(net_9985), .Z(net_12809) );
CLKBUF_X2 inst_13618 ( .A(net_13465), .Z(net_13466) );
INV_X4 inst_5192 ( .A(net_2846), .ZN(net_2845) );
CLKBUF_X2 inst_11566 ( .A(net_10516), .Z(net_11414) );
CLKBUF_X2 inst_11400 ( .A(net_11247), .Z(net_11248) );
CLKBUF_X2 inst_17501 ( .A(net_17348), .Z(net_17349) );
CLKBUF_X2 inst_12350 ( .A(net_12038), .Z(net_12198) );
CLKBUF_X2 inst_15406 ( .A(net_12946), .Z(net_15254) );
NAND4_X2 inst_3761 ( .ZN(net_4260), .A1(net_3824), .A2(net_3823), .A3(net_3822), .A4(net_3821) );
INV_X4 inst_5089 ( .ZN(net_5710), .A(net_5686) );
INV_X4 inst_5654 ( .A(net_6323), .ZN(net_644) );
CLKBUF_X2 inst_10138 ( .A(net_9519), .Z(net_9986) );
SDFF_X2 inst_853 ( .SI(net_8633), .Q(net_8633), .D(net_3977), .SE(net_3885), .CK(net_13319) );
INV_X4 inst_5864 ( .A(net_8923), .ZN(net_2612) );
SDFF_X2 inst_657 ( .Q(net_8430), .D(net_8430), .SI(net_3963), .SE(net_3934), .CK(net_10916) );
NAND2_X2 inst_4550 ( .A1(net_3369), .A2(net_3315), .ZN(net_3313) );
CLKBUF_X2 inst_12803 ( .A(net_12650), .Z(net_12651) );
SDFFS_X2 inst_2098 ( .Q(net_7526), .D(net_7526), .SI(net_1868), .SE(net_1136), .CK(net_16242), .SN(x6501) );
CLKBUF_X2 inst_12465 ( .A(net_12312), .Z(net_12313) );
SDFF_X2 inst_1921 ( .D(net_7284), .SI(net_6901), .Q(net_6901), .SE(net_6284), .CK(net_16167) );
CLKBUF_X2 inst_17467 ( .A(net_17314), .Z(net_17315) );
CLKBUF_X2 inst_12890 ( .A(net_12737), .Z(net_12738) );
CLKBUF_X2 inst_13890 ( .A(net_13119), .Z(net_13738) );
DFFR_X2 inst_6977 ( .QN(net_5974), .D(net_5904), .CK(net_11557), .RN(x6501) );
NAND2_X2 inst_4293 ( .A1(net_7130), .ZN(net_5167), .A2(net_5166) );
CLKBUF_X2 inst_13996 ( .A(net_13843), .Z(net_13844) );
CLKBUF_X2 inst_14783 ( .A(net_11629), .Z(net_14631) );
CLKBUF_X2 inst_10357 ( .A(net_9934), .Z(net_10205) );
CLKBUF_X2 inst_14285 ( .A(net_11433), .Z(net_14133) );
SDFFR_X2 inst_2638 ( .Q(net_7370), .D(net_7370), .SE(net_1136), .CK(net_18600), .RN(x6501), .SI(x4821) );
AOI222_X1 inst_8676 ( .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3335), .C1(net_3334), .A2(net_3172), .B1(net_3107) );
NOR4_X2 inst_3235 ( .ZN(net_1853), .A4(net_1573), .A2(net_946), .A1(net_929), .A3(net_925) );
CLKBUF_X2 inst_14019 ( .A(net_13866), .Z(net_13867) );
AOI222_X1 inst_8672 ( .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3545), .C1(net_3544), .A2(net_3235), .B1(net_3142) );
CLKBUF_X2 inst_14680 ( .A(net_11909), .Z(net_14528) );
CLKBUF_X2 inst_12786 ( .A(net_12633), .Z(net_12634) );
CLKBUF_X2 inst_9421 ( .A(net_9170), .Z(net_9269) );
AOI221_X4 inst_8711 ( .C1(net_8209), .B1(net_7699), .C2(net_6099), .ZN(net_6045), .B2(net_4399), .A(net_4289) );
AOI22_X2 inst_8125 ( .B1(net_8184), .A1(net_7674), .B2(net_6099), .A2(net_4399), .ZN(net_4024) );
SDFF_X2 inst_892 ( .Q(net_8578), .D(net_8578), .SI(net_3963), .SE(net_3878), .CK(net_12330) );
CLKBUF_X2 inst_17175 ( .A(net_17022), .Z(net_17023) );
NAND2_X2 inst_4100 ( .ZN(net_5433), .A1(net_5243), .A2(net_5014) );
CLKBUF_X2 inst_16053 ( .A(net_15900), .Z(net_15901) );
CLKBUF_X2 inst_17560 ( .A(net_17407), .Z(net_17408) );
SDFF_X2 inst_1803 ( .D(net_7295), .SI(net_6952), .Q(net_6952), .SE(net_6281), .CK(net_15424) );
DFFR_X2 inst_6987 ( .QN(net_5962), .D(net_5900), .CK(net_11494), .RN(x6501) );
OR2_X4 inst_2814 ( .ZN(net_5465), .A2(net_5461), .A1(net_4315) );
SDFF_X2 inst_936 ( .SI(net_7314), .Q(net_6655), .D(net_6655), .SE(net_3126), .CK(net_9960) );
CLKBUF_X2 inst_9819 ( .A(net_9666), .Z(net_9667) );
NAND4_X2 inst_3809 ( .ZN(net_3617), .A1(net_3451), .A2(net_3450), .A3(net_3449), .A4(net_3448) );
CLKBUF_X2 inst_14957 ( .A(net_14804), .Z(net_14805) );
CLKBUF_X2 inst_11368 ( .A(net_11215), .Z(net_11216) );
CLKBUF_X2 inst_14896 ( .A(net_14743), .Z(net_14744) );
CLKBUF_X2 inst_10315 ( .A(net_10162), .Z(net_10163) );
INV_X32 inst_6171 ( .ZN(net_5247), .A(net_4813) );
CLKBUF_X2 inst_14236 ( .A(net_14083), .Z(net_14084) );
CLKBUF_X2 inst_15300 ( .A(net_13720), .Z(net_15148) );
DFFS_X2 inst_6865 ( .QN(net_8971), .D(net_5281), .CK(net_17620), .SN(x6501) );
CLKBUF_X2 inst_12948 ( .A(net_11909), .Z(net_12796) );
NAND4_X2 inst_3780 ( .ZN(net_4241), .A1(net_3704), .A2(net_3703), .A3(net_3702), .A4(net_3701) );
SDFFR_X1 inst_2647 ( .D(net_6770), .SE(net_4506), .CK(net_9242), .RN(x6501), .SI(x1778), .Q(x1778) );
CLKBUF_X2 inst_11305 ( .A(net_9533), .Z(net_11153) );
CLKBUF_X2 inst_18938 ( .A(net_18785), .Z(net_18786) );
INV_X2 inst_6576 ( .A(net_8949), .ZN(net_607) );
CLKBUF_X2 inst_19090 ( .A(net_18937), .Z(net_18938) );
CLKBUF_X2 inst_15464 ( .A(net_11319), .Z(net_15312) );
SDFFR_X1 inst_2710 ( .SI(net_6815), .Q(net_6815), .D(net_6812), .SE(net_6267), .CK(net_11788), .RN(x6501) );
INV_X4 inst_5629 ( .A(net_7525), .ZN(net_1501) );
CLKBUF_X2 inst_11959 ( .A(net_11806), .Z(net_11807) );
SDFF_X2 inst_1058 ( .D(net_7313), .SI(net_6621), .Q(net_6621), .SE(net_3123), .CK(net_12014) );
CLKBUF_X2 inst_12639 ( .A(net_12486), .Z(net_12487) );
NOR2_X2 inst_3360 ( .ZN(net_5565), .A2(net_5388), .A1(net_5387) );
DFF_X1 inst_6821 ( .QN(net_8235), .D(net_4446), .CK(net_17200) );
CLKBUF_X2 inst_16441 ( .A(net_11176), .Z(net_16289) );
MUX2_X2 inst_4984 ( .A(net_9041), .Z(net_3975), .B(net_3224), .S(net_622) );
CLKBUF_X2 inst_18539 ( .A(net_12123), .Z(net_18387) );
CLKBUF_X2 inst_18206 ( .A(net_17596), .Z(net_18054) );
SDFF_X2 inst_1788 ( .SI(net_8068), .Q(net_8068), .D(net_2717), .SE(net_2508), .CK(net_16464) );
CLKBUF_X2 inst_14098 ( .A(net_13945), .Z(net_13946) );
SDFF_X2 inst_1272 ( .Q(net_8083), .D(net_8083), .SE(net_2707), .SI(net_2659), .CK(net_15300) );
CLKBUF_X2 inst_17780 ( .A(net_11321), .Z(net_17628) );
NAND2_X2 inst_4182 ( .ZN(net_5321), .A2(net_5188), .A1(net_5072) );
CLKBUF_X2 inst_14566 ( .A(net_14413), .Z(net_14414) );
OR2_X4 inst_2852 ( .ZN(net_6086), .A1(net_772), .A2(net_476) );
DFF_X1 inst_6751 ( .Q(net_6761), .D(net_5615), .CK(net_10494) );
CLKBUF_X2 inst_17008 ( .A(net_16855), .Z(net_16856) );
CLKBUF_X2 inst_18458 ( .A(net_18305), .Z(net_18306) );
NAND3_X2 inst_3973 ( .A3(net_9008), .A2(net_6119), .ZN(net_2423), .A1(net_1821) );
SDFF_X2 inst_433 ( .Q(net_8761), .D(net_8761), .SE(net_3982), .SI(net_3957), .CK(net_13286) );
CLKBUF_X2 inst_13771 ( .A(net_13618), .Z(net_13619) );
MUX2_X2 inst_4939 ( .S(net_2963), .Z(net_2784), .A(net_2311), .B(net_553) );
CLKBUF_X2 inst_11817 ( .A(net_9470), .Z(net_11665) );
CLKBUF_X2 inst_13249 ( .A(net_11249), .Z(net_13097) );
CLKBUF_X2 inst_18925 ( .A(net_17366), .Z(net_18773) );
CLKBUF_X2 inst_17605 ( .A(net_16719), .Z(net_17453) );
CLKBUF_X2 inst_18454 ( .A(net_18301), .Z(net_18302) );
INV_X2 inst_6417 ( .ZN(net_810), .A(net_809) );
CLKBUF_X2 inst_11312 ( .A(net_11159), .Z(net_11160) );
CLKBUF_X2 inst_13772 ( .A(net_13619), .Z(net_13620) );
AOI21_X2 inst_8984 ( .ZN(net_1890), .B2(net_1883), .A(net_1812), .B1(net_1140) );
CLKBUF_X2 inst_16411 ( .A(net_13695), .Z(net_16259) );
CLKBUF_X2 inst_11955 ( .A(net_11802), .Z(net_11803) );
AOI222_X1 inst_8638 ( .C2(net_5832), .A2(net_5830), .B2(net_5824), .ZN(net_3988), .A1(net_3541), .B1(net_2134), .C1(x2856) );
CLKBUF_X2 inst_9269 ( .A(net_9093), .Z(net_9117) );
INV_X4 inst_5781 ( .A(net_7205), .ZN(net_2953) );
CLKBUF_X2 inst_13476 ( .A(net_11609), .Z(net_13324) );
CLKBUF_X2 inst_14733 ( .A(net_14580), .Z(net_14581) );
DFFR_X2 inst_7151 ( .QN(net_6400), .D(net_2823), .CK(net_17935), .RN(x6501) );
CLKBUF_X2 inst_15325 ( .A(net_12298), .Z(net_15173) );
CLKBUF_X2 inst_17564 ( .A(net_17411), .Z(net_17412) );
SDFF_X2 inst_1475 ( .SI(net_7270), .Q(net_7127), .D(net_7127), .SE(net_6279), .CK(net_16841) );
CLKBUF_X2 inst_15960 ( .A(net_15807), .Z(net_15808) );
SDFF_X2 inst_1637 ( .Q(net_8152), .D(net_8152), .SI(net_2708), .SE(net_2538), .CK(net_15513) );
SDFF_X2 inst_1352 ( .SI(net_7843), .Q(net_7843), .D(net_2655), .SE(net_2558), .CK(net_15464) );
CLKBUF_X2 inst_17079 ( .A(net_9194), .Z(net_16927) );
CLKBUF_X2 inst_12338 ( .A(net_12185), .Z(net_12186) );
SDFFR_X2 inst_2261 ( .D(net_7392), .SE(net_2801), .SI(net_201), .Q(net_201), .CK(net_14979), .RN(x6501) );
CLKBUF_X2 inst_9955 ( .A(net_9073), .Z(net_9803) );
CLKBUF_X2 inst_18374 ( .A(net_13382), .Z(net_18222) );
CLKBUF_X2 inst_14524 ( .A(net_14371), .Z(net_14372) );
NOR2_X2 inst_3390 ( .A2(net_4553), .ZN(net_4474), .A1(net_1688) );
AND2_X4 inst_9076 ( .ZN(net_3215), .A2(net_3176), .A1(net_3157) );
CLKBUF_X2 inst_15742 ( .A(net_9328), .Z(net_15590) );
CLKBUF_X2 inst_16945 ( .A(net_16792), .Z(net_16793) );
OAI22_X2 inst_2930 ( .A2(net_2650), .B2(net_2649), .ZN(net_2485), .A1(net_1044), .B1(net_768) );
AOI22_X2 inst_8178 ( .B1(net_8752), .A1(net_8382), .A2(net_3867), .B2(net_3866), .ZN(net_3853) );
INV_X4 inst_5683 ( .ZN(net_2742), .A(net_277) );
NAND2_X2 inst_4790 ( .ZN(net_4380), .A2(net_1504), .A1(net_1355) );
NAND2_X2 inst_4307 ( .A1(net_7054), .A2(net_5162), .ZN(net_5150) );
CLKBUF_X2 inst_9851 ( .A(net_9698), .Z(net_9699) );
CLKBUF_X2 inst_18082 ( .A(net_11822), .Z(net_17930) );
OAI211_X2 inst_3192 ( .C1(net_7212), .ZN(net_3164), .A(net_3163), .B(net_1728), .C2(net_1727) );
MUX2_X2 inst_5006 ( .A(net_9046), .Z(net_3951), .B(net_3921), .S(net_622) );
AND4_X4 inst_9026 ( .ZN(net_4968), .A4(net_4719), .A1(net_4575), .A2(net_4536), .A3(net_4480) );
CLKBUF_X2 inst_18485 ( .A(net_18332), .Z(net_18333) );
CLKBUF_X2 inst_9780 ( .A(net_9627), .Z(net_9628) );
CLKBUF_X2 inst_19078 ( .A(net_18925), .Z(net_18926) );
CLKBUF_X2 inst_13585 ( .A(net_13432), .Z(net_13433) );
CLKBUF_X2 inst_11129 ( .A(net_10722), .Z(net_10977) );
NAND2_X2 inst_4246 ( .A1(net_7026), .A2(net_5249), .ZN(net_5214) );
AND2_X4 inst_9146 ( .A1(net_7523), .A2(net_6323), .ZN(net_1089) );
NAND3_X2 inst_3904 ( .ZN(net_5634), .A1(net_5563), .A3(net_5497), .A2(net_5378) );
CLKBUF_X2 inst_10634 ( .A(net_10481), .Z(net_10482) );
INV_X2 inst_6333 ( .ZN(net_3004), .A(net_2964) );
INV_X4 inst_5649 ( .A(net_7384), .ZN(net_945) );
SDFF_X2 inst_1393 ( .SI(net_7727), .Q(net_7727), .D(net_2749), .SE(net_2559), .CK(net_13782) );
INV_X2 inst_6276 ( .ZN(net_4319), .A(net_4318) );
NOR2_X2 inst_3519 ( .ZN(net_1751), .A1(net_1750), .A2(net_1749) );
NAND2_X2 inst_4075 ( .A2(net_6767), .A1(net_5835), .ZN(net_5771) );
CLKBUF_X2 inst_13402 ( .A(net_13249), .Z(net_13250) );
CLKBUF_X2 inst_16191 ( .A(net_16038), .Z(net_16039) );
CLKBUF_X2 inst_17948 ( .A(net_15949), .Z(net_17796) );
CLKBUF_X2 inst_15720 ( .A(net_15567), .Z(net_15568) );
CLKBUF_X2 inst_16576 ( .A(net_16423), .Z(net_16424) );
INV_X4 inst_5153 ( .ZN(net_3211), .A(net_3175) );
INV_X4 inst_5731 ( .A(net_8930), .ZN(net_4551) );
CLKBUF_X2 inst_14264 ( .A(net_14111), .Z(net_14112) );
CLKBUF_X2 inst_15913 ( .A(net_15760), .Z(net_15761) );
AOI222_X1 inst_8631 ( .A2(net_6452), .A1(net_5654), .C2(net_5595), .B2(net_4881), .ZN(net_4706), .C1(net_334), .B1(net_252) );
CLKBUF_X2 inst_13118 ( .A(net_12965), .Z(net_12966) );
CLKBUF_X2 inst_14446 ( .A(net_12429), .Z(net_14294) );
CLKBUF_X2 inst_18610 ( .A(net_15781), .Z(net_18458) );
NAND2_X2 inst_4791 ( .ZN(net_3262), .A2(net_1503), .A1(net_501) );
INV_X2 inst_6459 ( .A(net_7569), .ZN(net_3130) );
AOI22_X2 inst_8007 ( .B1(net_8181), .A1(net_7671), .B2(net_6099), .A2(net_4399), .ZN(net_4127) );
CLKBUF_X2 inst_15866 ( .A(net_15713), .Z(net_15714) );
OAI22_X2 inst_2937 ( .ZN(net_2044), .A1(net_2043), .B1(net_1833), .A2(net_1794), .B2(net_1136) );
DFFR_X2 inst_7244 ( .QN(net_7232), .D(net_2065), .CK(net_17783), .RN(x6501) );
CLKBUF_X2 inst_17124 ( .A(net_16971), .Z(net_16972) );
SDFF_X2 inst_687 ( .Q(net_8860), .D(net_8860), .SI(net_3937), .SE(net_3936), .CK(net_12442) );
AOI22_X2 inst_7864 ( .B2(net_4881), .A2(net_4809), .ZN(net_4577), .A1(net_348), .B1(net_254) );
SDFFR_X2 inst_2319 ( .SE(net_2260), .Q(net_381), .D(net_381), .CK(net_11399), .RN(x6501), .SI(x1281) );
DFFR_X2 inst_7091 ( .QN(net_8291), .D(net_3553), .CK(net_12060), .RN(x6501) );
INV_X4 inst_5519 ( .A(net_1756), .ZN(net_674) );
SDFFR_X2 inst_2225 ( .Q(net_7470), .D(net_7470), .SE(net_2863), .CK(net_12182), .SI(x13433), .RN(x6501) );
AOI22_X2 inst_7927 ( .B1(net_8112), .A1(net_7874), .A2(net_6098), .ZN(net_4197), .B2(net_4190) );
CLKBUF_X2 inst_16523 ( .A(net_16370), .Z(net_16371) );
CLKBUF_X2 inst_13805 ( .A(net_13652), .Z(net_13653) );
CLKBUF_X2 inst_17889 ( .A(net_17263), .Z(net_17737) );
CLKBUF_X2 inst_17428 ( .A(net_12753), .Z(net_17276) );
NAND2_X2 inst_4061 ( .ZN(net_5880), .A2(net_5768), .A1(net_3585) );
SDFFR_X2 inst_2513 ( .D(net_7366), .SI(net_2501), .SE(net_2225), .QN(net_339), .CK(net_16102), .RN(x6501) );
SDFFR_X2 inst_2254 ( .D(net_7366), .SI(net_2800), .SE(net_2442), .QN(net_266), .CK(net_16137), .RN(x6501) );
CLKBUF_X2 inst_14690 ( .A(net_9206), .Z(net_14538) );
AOI22_X2 inst_7775 ( .B1(net_6965), .A1(net_6925), .A2(net_5443), .B2(net_5442), .ZN(net_5303) );
CLKBUF_X2 inst_18844 ( .A(net_18691), .Z(net_18692) );
INV_X2 inst_6255 ( .ZN(net_4734), .A(net_4690) );
CLKBUF_X2 inst_10111 ( .A(net_9958), .Z(net_9959) );
CLKBUF_X2 inst_9255 ( .A(net_9102), .Z(net_9103) );
CLKBUF_X2 inst_16531 ( .A(net_16378), .Z(net_16379) );
CLKBUF_X2 inst_10922 ( .A(net_9954), .Z(net_10770) );
CLKBUF_X2 inst_12519 ( .A(net_12366), .Z(net_12367) );
CLKBUF_X2 inst_15479 ( .A(net_15326), .Z(net_15327) );
CLKBUF_X2 inst_16640 ( .A(net_16487), .Z(net_16488) );
CLKBUF_X2 inst_11755 ( .A(net_11602), .Z(net_11603) );
SDFF_X2 inst_354 ( .Q(net_8774), .D(net_8774), .SE(net_3982), .SI(net_3976), .CK(net_12645) );
CLKBUF_X2 inst_13794 ( .A(net_13641), .Z(net_13642) );
SDFF_X2 inst_1145 ( .SI(net_7325), .Q(net_6600), .D(net_6600), .SE(net_3069), .CK(net_9122) );
INV_X2 inst_6235 ( .ZN(net_5475), .A(net_5286) );
CLKBUF_X2 inst_12859 ( .A(net_12706), .Z(net_12707) );
CLKBUF_X2 inst_15380 ( .A(net_15227), .Z(net_15228) );
CLKBUF_X2 inst_15981 ( .A(net_15828), .Z(net_15829) );
CLKBUF_X2 inst_18545 ( .A(net_18392), .Z(net_18393) );
CLKBUF_X2 inst_14804 ( .A(net_9294), .Z(net_14652) );
CLKBUF_X1 inst_7731 ( .A(x192486), .Z(x1032) );
CLKBUF_X2 inst_16006 ( .A(net_11668), .Z(net_15854) );
CLKBUF_X2 inst_16521 ( .A(net_16368), .Z(net_16369) );
AOI22_X2 inst_8414 ( .B1(net_8565), .A1(net_8454), .A2(net_6263), .B2(net_6262), .ZN(net_3638) );
SDFF_X2 inst_1717 ( .Q(net_8004), .D(net_8004), .SI(net_2715), .SE(net_2542), .CK(net_14159) );
CLKBUF_X2 inst_18359 ( .A(net_18206), .Z(net_18207) );
CLKBUF_X2 inst_15206 ( .A(net_15053), .Z(net_15054) );
OR2_X2 inst_2901 ( .A2(net_7306), .A1(net_7305), .ZN(net_809) );
INV_X4 inst_6080 ( .A(net_7586), .ZN(net_491) );
SDFF_X2 inst_718 ( .SI(net_8644), .Q(net_8644), .D(net_3959), .SE(net_3885), .CK(net_13188) );
CLKBUF_X2 inst_17488 ( .A(net_17259), .Z(net_17336) );
CLKBUF_X2 inst_17707 ( .A(net_17554), .Z(net_17555) );
NAND2_X4 inst_4024 ( .ZN(net_6195), .A2(net_3362), .A1(net_3308) );
CLKBUF_X2 inst_18254 ( .A(net_18101), .Z(net_18102) );
DFFR_X2 inst_7362 ( .Q(net_7320), .CK(net_11360), .D(x13093), .RN(x6501) );
AOI22_X2 inst_8100 ( .B1(net_8212), .A1(net_7702), .B2(net_6099), .A2(net_4399), .ZN(net_4048) );
AND2_X2 inst_9166 ( .ZN(net_2809), .A2(net_2554), .A1(net_1159) );
INV_X4 inst_5585 ( .A(net_7571), .ZN(net_595) );
AOI22_X2 inst_8350 ( .B1(net_8738), .A1(net_8516), .B2(net_4350), .A2(net_4349), .ZN(net_3698) );
CLKBUF_X2 inst_17827 ( .A(net_17674), .Z(net_17675) );
SDFFR_X2 inst_2147 ( .QN(net_8260), .D(net_2997), .SE(net_2996), .SI(net_1231), .CK(net_18461), .RN(x6501) );
CLKBUF_X2 inst_13171 ( .A(net_13018), .Z(net_13019) );
SDFFS_X2 inst_2091 ( .SI(net_6835), .Q(net_6835), .SE(net_2146), .D(net_1218), .CK(net_18673), .SN(x6501) );
CLKBUF_X2 inst_19135 ( .A(net_18982), .Z(net_18983) );
CLKBUF_X2 inst_18423 ( .A(net_18270), .Z(net_18271) );
CLKBUF_X2 inst_10733 ( .A(net_9063), .Z(net_10581) );
CLKBUF_X2 inst_12247 ( .A(net_12094), .Z(net_12095) );
AOI22_X2 inst_8066 ( .B1(net_8106), .A1(net_7766), .B2(net_6108), .A2(net_6096), .ZN(net_4077) );
INV_X4 inst_5863 ( .A(net_6823), .ZN(net_990) );
CLKBUF_X2 inst_16783 ( .A(net_16630), .Z(net_16631) );
SDFF_X2 inst_500 ( .SI(net_8626), .Q(net_8626), .SE(net_3984), .D(net_3976), .CK(net_10368) );
INV_X4 inst_5348 ( .A(net_3003), .ZN(net_1705) );
CLKBUF_X2 inst_14403 ( .A(net_14250), .Z(net_14251) );
SDFF_X2 inst_550 ( .Q(net_8695), .D(net_8695), .SI(net_3953), .SE(net_3935), .CK(net_10270) );
DFF_X1 inst_6758 ( .Q(net_7539), .D(net_4613), .CK(net_9739) );
CLKBUF_X2 inst_16270 ( .A(net_16117), .Z(net_16118) );
CLKBUF_X2 inst_17213 ( .A(net_10183), .Z(net_17061) );
INV_X4 inst_5913 ( .A(net_7425), .ZN(net_3330) );
CLKBUF_X2 inst_11972 ( .A(net_11819), .Z(net_11820) );
CLKBUF_X2 inst_13610 ( .A(net_11055), .Z(net_13458) );
AOI22_X2 inst_8311 ( .B1(net_8881), .A1(net_8326), .B2(net_6252), .A2(net_4345), .ZN(net_3734) );
CLKBUF_X2 inst_17761 ( .A(net_17608), .Z(net_17609) );
AOI222_X1 inst_8702 ( .A1(net_5031), .B2(net_5028), .C2(net_5027), .ZN(net_2792), .A2(net_2791), .B1(net_2790), .C1(net_1536) );
CLKBUF_X2 inst_15417 ( .A(net_15264), .Z(net_15265) );
INV_X4 inst_5471 ( .ZN(net_874), .A(net_747) );
SDFFR_X1 inst_2661 ( .D(net_6783), .SE(net_4506), .CK(net_11408), .RN(x6501), .SI(x1340), .Q(x1340) );
AOI22_X2 inst_8237 ( .B1(net_8705), .A1(net_8483), .B2(net_4350), .A2(net_4349), .ZN(net_3800) );
INV_X4 inst_6034 ( .A(net_7433), .ZN(net_3990) );
NOR2_X2 inst_3548 ( .ZN(net_1443), .A2(net_1442), .A1(net_1153) );
CLKBUF_X2 inst_15246 ( .A(net_15093), .Z(net_15094) );
SDFF_X2 inst_594 ( .SI(net_8386), .Q(net_8386), .D(net_3973), .SE(net_3969), .CK(net_10841) );
CLKBUF_X2 inst_13848 ( .A(net_13695), .Z(net_13696) );
NAND2_X2 inst_4435 ( .A1(net_6872), .A2(net_5016), .ZN(net_4992) );
SDFFR_X2 inst_2175 ( .QN(net_9009), .SE(net_2960), .SI(net_2959), .D(net_915), .CK(net_11198), .RN(x6501) );
SDFF_X2 inst_1632 ( .Q(net_8177), .D(net_8177), .SI(net_2716), .SE(net_2538), .CK(net_17065) );
NAND2_X2 inst_4241 ( .A1(net_6903), .A2(net_5247), .ZN(net_5219) );
SDFF_X2 inst_925 ( .SI(net_8732), .Q(net_8732), .SE(net_6195), .D(net_3953), .CK(net_10211) );
SDFFR_X2 inst_2193 ( .SE(net_6752), .Q(net_6752), .SI(net_2933), .D(net_2897), .CK(net_9112), .RN(x6501) );
CLKBUF_X2 inst_10302 ( .A(net_9085), .Z(net_10150) );
AOI221_X4 inst_8734 ( .B1(net_8740), .C1(net_8518), .B2(net_4350), .C2(net_4349), .ZN(net_4332), .A(net_4238) );
CLKBUF_X2 inst_9793 ( .A(net_9187), .Z(net_9641) );
INV_X4 inst_6147 ( .A(net_6809), .ZN(net_6142) );
AOI21_X2 inst_8999 ( .ZN(net_1275), .A(net_1274), .B1(net_1273), .B2(net_841) );
SDFF_X2 inst_881 ( .Q(net_8560), .D(net_8560), .SI(net_3938), .SE(net_3878), .CK(net_12409) );
SDFF_X2 inst_1536 ( .Q(net_7988), .D(net_7988), .SI(net_2574), .SE(net_2542), .CK(net_15593) );
NAND3_X4 inst_3876 ( .ZN(net_2459), .A1(net_2299), .A3(net_2088), .A2(net_1694) );
CLKBUF_X2 inst_11300 ( .A(net_11147), .Z(net_11148) );
NAND4_X2 inst_3848 ( .ZN(net_1719), .A4(net_1244), .A2(net_1022), .A1(net_1000), .A3(net_963) );
DFFR_X2 inst_7001 ( .D(net_5879), .CK(net_11440), .RN(x6501), .Q(x2594) );
CLKBUF_X2 inst_12175 ( .A(net_9386), .Z(net_12023) );
CLKBUF_X2 inst_19034 ( .A(net_18881), .Z(net_18882) );
NAND4_X2 inst_3706 ( .A4(net_6232), .A1(net_6231), .ZN(net_4431), .A2(net_3726), .A3(net_3725) );
CLKBUF_X2 inst_13979 ( .A(net_13826), .Z(net_13827) );
CLKBUF_X2 inst_9219 ( .A(net_9066), .Z(net_9067) );
XNOR2_X2 inst_247 ( .A(net_2726), .B(net_2679), .ZN(net_1204) );
SDFF_X2 inst_403 ( .SI(net_8316), .Q(net_8316), .SE(net_3978), .D(net_3974), .CK(net_12289) );
INV_X4 inst_6089 ( .A(net_7165), .ZN(net_864) );
DFFR_X2 inst_7066 ( .QN(net_7419), .D(net_4200), .CK(net_12310), .RN(x6501) );
CLKBUF_X2 inst_17727 ( .A(net_17574), .Z(net_17575) );
CLKBUF_X2 inst_15969 ( .A(net_15816), .Z(net_15817) );
CLKBUF_X2 inst_15883 ( .A(net_9127), .Z(net_15731) );
NOR2_X2 inst_3446 ( .ZN(net_3024), .A1(net_3023), .A2(net_2930) );
SDFFR_X1 inst_2728 ( .SI(net_9041), .Q(net_9041), .D(net_7470), .SE(net_3208), .CK(net_12219), .RN(x6501) );
CLKBUF_X2 inst_16559 ( .A(net_9428), .Z(net_16407) );
SDFF_X2 inst_1588 ( .Q(net_8014), .D(net_8014), .SI(net_2709), .SE(net_2545), .CK(net_15768) );
CLKBUF_X2 inst_18790 ( .A(net_18637), .Z(net_18638) );
CLKBUF_X2 inst_18310 ( .A(net_18157), .Z(net_18158) );
AOI22_X2 inst_8002 ( .A1(net_7943), .B1(net_7773), .A2(net_6092), .B2(net_6091), .ZN(net_4132) );
CLKBUF_X2 inst_14484 ( .A(net_14331), .Z(net_14332) );
CLKBUF_X2 inst_10996 ( .A(net_10843), .Z(net_10844) );
SDFFR_X2 inst_2516 ( .QN(net_6409), .SE(net_2218), .SI(net_2217), .D(net_1843), .CK(net_9611), .RN(x6501) );
CLKBUF_X2 inst_13901 ( .A(net_13748), .Z(net_13749) );
SDFF_X2 inst_1506 ( .SI(net_7866), .Q(net_7866), .D(net_2710), .SE(net_2558), .CK(net_14419) );
CLKBUF_X2 inst_9567 ( .A(net_9212), .Z(net_9415) );
CLKBUF_X2 inst_9494 ( .A(net_9341), .Z(net_9342) );
CLKBUF_X2 inst_15515 ( .A(net_15362), .Z(net_15363) );
NAND4_X2 inst_3785 ( .ZN(net_4236), .A1(net_3670), .A2(net_3669), .A3(net_3668), .A4(net_3667) );
INV_X4 inst_6058 ( .ZN(net_2546), .A(net_259) );
DFFR_X1 inst_7541 ( .Q(net_7654), .D(net_917), .CK(net_12708), .RN(x6501) );
CLKBUF_X2 inst_10455 ( .A(net_10302), .Z(net_10303) );
CLKBUF_X2 inst_16987 ( .A(net_16087), .Z(net_16835) );
CLKBUF_X2 inst_15800 ( .A(net_15647), .Z(net_15648) );
INV_X4 inst_5678 ( .A(net_7646), .ZN(net_738) );
DFFR_X1 inst_7454 ( .QN(net_8939), .D(net_4742), .CK(net_13742), .RN(x6501) );
SDFF_X2 inst_1361 ( .SI(net_7845), .Q(net_7845), .D(net_2659), .SE(net_2558), .CK(net_18562) );
NOR2_X2 inst_3401 ( .A2(net_6206), .ZN(net_4317), .A1(net_4316) );
CLKBUF_X2 inst_12949 ( .A(net_10651), .Z(net_12797) );
CLKBUF_X2 inst_13105 ( .A(net_12952), .Z(net_12953) );
CLKBUF_X2 inst_12688 ( .A(net_12535), .Z(net_12536) );
DFFR_X1 inst_7525 ( .Q(net_7661), .D(net_7657), .CK(net_12720), .RN(x6501) );
CLKBUF_X2 inst_11916 ( .A(net_11763), .Z(net_11764) );
CLKBUF_X2 inst_12439 ( .A(net_12286), .Z(net_12287) );
SDFFR_X2 inst_2208 ( .Q(net_7463), .D(net_7463), .SE(net_2863), .CK(net_10635), .SI(x13488), .RN(x6501) );
NAND2_X2 inst_4463 ( .ZN(net_4785), .A2(net_4783), .A1(x1215) );
CLKBUF_X2 inst_18410 ( .A(net_10568), .Z(net_18258) );
INV_X4 inst_5598 ( .A(net_6423), .ZN(net_1829) );
AOI221_X2 inst_8789 ( .C2(net_5609), .ZN(net_4966), .B2(net_4965), .A(net_4695), .B1(net_2737), .C1(net_357) );
CLKBUF_X2 inst_10698 ( .A(net_10545), .Z(net_10546) );
AOI21_X2 inst_8975 ( .ZN(net_2539), .B2(net_2204), .A(net_2103), .B1(net_1261) );
AOI22_X2 inst_7873 ( .A2(net_6438), .A1(net_5654), .B2(net_4881), .ZN(net_4568), .B1(net_238) );
SDFFR_X2 inst_2174 ( .QN(net_7599), .SE(net_3144), .D(net_3127), .SI(net_1093), .CK(net_13500), .RN(x6501) );
DFF_X1 inst_6721 ( .Q(net_6767), .D(net_5648), .CK(net_9268) );
CLKBUF_X2 inst_10779 ( .A(net_10617), .Z(net_10627) );
CLKBUF_X2 inst_13089 ( .A(net_12374), .Z(net_12937) );
XOR2_X2 inst_14 ( .Z(net_1490), .A(net_1489), .B(net_1343) );
AOI22_X2 inst_7886 ( .B1(net_8997), .A2(net_5538), .B2(net_5456), .ZN(net_4545), .A1(net_426) );
CLKBUF_X2 inst_9366 ( .A(net_9213), .Z(net_9214) );
DFFR_X2 inst_7172 ( .QN(net_6169), .D(net_2509), .CK(net_11217), .RN(x6501) );
CLKBUF_X2 inst_15774 ( .A(net_15621), .Z(net_15622) );
CLKBUF_X2 inst_15085 ( .A(net_12414), .Z(net_14933) );
SDFFR_X2 inst_2325 ( .SE(net_2260), .Q(net_374), .D(net_374), .CK(net_11466), .RN(x6501), .SI(x1532) );
CLKBUF_X2 inst_12068 ( .A(net_11915), .Z(net_11916) );
CLKBUF_X2 inst_12354 ( .A(net_12201), .Z(net_12202) );
SDFF_X2 inst_1074 ( .D(net_7323), .SI(net_6499), .Q(net_6499), .SE(net_3071), .CK(net_11351) );
AOI22_X2 inst_7983 ( .B1(net_8061), .A1(net_7857), .B2(net_6107), .A2(net_4400), .ZN(net_4148) );
DFFR_X1 inst_7375 ( .QN(net_5943), .D(net_5886), .CK(net_9402), .RN(x6501) );
CLKBUF_X2 inst_10149 ( .A(net_9259), .Z(net_9997) );
CLKBUF_X2 inst_14944 ( .A(net_9784), .Z(net_14792) );
SDFF_X2 inst_1602 ( .Q(net_8138), .D(net_8138), .SI(net_2710), .SE(net_2541), .CK(net_16485) );
CLKBUF_X2 inst_9883 ( .A(net_9730), .Z(net_9731) );
CLKBUF_X2 inst_11100 ( .A(net_10129), .Z(net_10948) );
SDFF_X2 inst_969 ( .SI(net_7330), .Q(net_6737), .D(net_6737), .SE(net_3124), .CK(net_9103) );
CLKBUF_X2 inst_14569 ( .A(net_14416), .Z(net_14417) );
CLKBUF_X2 inst_18465 ( .A(net_18312), .Z(net_18313) );
INV_X2 inst_6463 ( .A(net_7423), .ZN(net_578) );
AOI22_X2 inst_8567 ( .ZN(net_2173), .A2(net_2172), .B1(net_2133), .A1(net_2071), .B2(net_1820) );
CLKBUF_X2 inst_13081 ( .A(net_11376), .Z(net_12929) );
SDFFR_X2 inst_2528 ( .D(net_7368), .SE(net_2387), .SI(net_283), .Q(net_283), .CK(net_13669), .RN(x6501) );
CLKBUF_X2 inst_12487 ( .A(net_11483), .Z(net_12335) );
CLKBUF_X2 inst_17534 ( .A(net_17381), .Z(net_17382) );
MUX2_X2 inst_4917 ( .B(net_6321), .Z(net_5524), .A(net_5523), .S(net_5522) );
CLKBUF_X2 inst_9749 ( .A(net_9596), .Z(net_9597) );
DFFR_X2 inst_7049 ( .QN(net_7497), .D(net_4724), .CK(net_17250), .RN(x6501) );
NAND2_X2 inst_4227 ( .A1(net_6897), .A2(net_5247), .ZN(net_5233) );
DFF_X1 inst_6840 ( .Q(net_6430), .D(net_3607), .CK(net_17977) );
CLKBUF_X2 inst_9800 ( .A(net_9647), .Z(net_9648) );
CLKBUF_X2 inst_16599 ( .A(net_10253), .Z(net_16447) );
CLKBUF_X2 inst_10824 ( .A(net_10671), .Z(net_10672) );
CLKBUF_X2 inst_18478 ( .A(net_15469), .Z(net_18326) );
CLKBUF_X2 inst_12290 ( .A(net_9320), .Z(net_12138) );
SDFFR_X2 inst_2343 ( .SI(net_7380), .D(net_2735), .SE(net_2723), .QN(net_161), .CK(net_17818), .RN(x6501) );
SDFFR_X2 inst_2538 ( .QN(net_6377), .SE(net_2147), .D(net_2144), .SI(net_1953), .CK(net_18147), .RN(x6501) );
CLKBUF_X2 inst_11500 ( .A(net_11347), .Z(net_11348) );
INV_X4 inst_5708 ( .A(net_8942), .ZN(net_1028) );
CLKBUF_X2 inst_12303 ( .A(net_9794), .Z(net_12151) );
CLKBUF_X2 inst_16980 ( .A(net_16827), .Z(net_16828) );
CLKBUF_X2 inst_12427 ( .A(net_12274), .Z(net_12275) );
CLKBUF_X2 inst_11929 ( .A(net_10207), .Z(net_11777) );
CLKBUF_X2 inst_15599 ( .A(net_15446), .Z(net_15447) );
CLKBUF_X2 inst_12584 ( .A(net_12431), .Z(net_12432) );
MUX2_X2 inst_4945 ( .S(net_3354), .Z(net_2521), .B(net_2520), .A(net_2109) );
INV_X4 inst_5169 ( .ZN(net_5912), .A(net_5832) );
AOI221_X2 inst_8782 ( .B1(net_7189), .C2(net_6187), .B2(net_5655), .ZN(net_5256), .A(net_4932), .C1(net_190) );
CLKBUF_X2 inst_15497 ( .A(net_13374), .Z(net_15345) );
CLKBUF_X2 inst_9982 ( .A(net_9829), .Z(net_9830) );
CLKBUF_X2 inst_17519 ( .A(net_17366), .Z(net_17367) );
CLKBUF_X2 inst_10970 ( .A(net_9906), .Z(net_10818) );
CLKBUF_X2 inst_13908 ( .A(net_10562), .Z(net_13756) );
SDFF_X2 inst_1089 ( .D(net_7310), .SI(net_6519), .Q(net_6519), .SE(net_3071), .CK(net_11875) );
CLKBUF_X2 inst_9720 ( .A(net_9567), .Z(net_9568) );
CLKBUF_X2 inst_17198 ( .A(net_15396), .Z(net_17046) );
INV_X2 inst_6537 ( .A(net_7564), .ZN(net_3108) );
CLKBUF_X2 inst_10251 ( .A(net_10098), .Z(net_10099) );
INV_X2 inst_6430 ( .ZN(net_6215), .A(net_1039) );
CLKBUF_X2 inst_17586 ( .A(net_17433), .Z(net_17434) );
DFFS_X1 inst_6932 ( .D(net_6145), .CK(net_16353), .SN(x6501), .Q(x871) );
INV_X4 inst_5367 ( .ZN(net_1135), .A(net_1134) );
AND2_X4 inst_9092 ( .ZN(net_2755), .A2(net_2381), .A1(net_2263) );
CLKBUF_X2 inst_12614 ( .A(net_9546), .Z(net_12462) );
CLKBUF_X2 inst_17127 ( .A(net_16974), .Z(net_16975) );
SDFF_X2 inst_2046 ( .SI(net_7805), .Q(net_7805), .D(net_2703), .SE(net_2459), .CK(net_13989) );
INV_X4 inst_6041 ( .A(net_7582), .ZN(net_749) );
CLKBUF_X2 inst_12021 ( .A(net_11357), .Z(net_11869) );
NAND2_X2 inst_4129 ( .ZN(net_5395), .A2(net_5224), .A1(net_5126) );
DFFR_X1 inst_7505 ( .D(net_1818), .Q(net_296), .CK(net_11187), .RN(x6501) );
CLKBUF_X2 inst_11632 ( .A(net_11479), .Z(net_11480) );
INV_X2 inst_6340 ( .ZN(net_2841), .A(net_2591) );
CLKBUF_X2 inst_18453 ( .A(net_18300), .Z(net_18301) );
CLKBUF_X2 inst_14176 ( .A(net_12317), .Z(net_14024) );
CLKBUF_X2 inst_16410 ( .A(net_16257), .Z(net_16258) );
CLKBUF_X2 inst_15953 ( .A(net_13485), .Z(net_15801) );
CLKBUF_X2 inst_14835 ( .A(net_12473), .Z(net_14683) );
CLKBUF_X2 inst_19121 ( .A(net_15798), .Z(net_18969) );
CLKBUF_X2 inst_13783 ( .A(net_13148), .Z(net_13631) );
CLKBUF_X2 inst_14224 ( .A(net_14071), .Z(net_14072) );
CLKBUF_X2 inst_15833 ( .A(net_13085), .Z(net_15681) );
INV_X2 inst_6533 ( .A(net_7565), .ZN(net_3133) );
CLKBUF_X2 inst_17510 ( .A(net_9936), .Z(net_17358) );
NOR2_X2 inst_3524 ( .ZN(net_6276), .A2(net_6123), .A1(net_1716) );
NAND2_X2 inst_4479 ( .A2(net_4624), .ZN(net_4504), .A1(net_1830) );
CLKBUF_X2 inst_12333 ( .A(net_12180), .Z(net_12181) );
CLKBUF_X2 inst_10882 ( .A(net_10191), .Z(net_10730) );
NAND2_X2 inst_4782 ( .ZN(net_1578), .A1(net_1577), .A2(net_1576) );
CLKBUF_X2 inst_15283 ( .A(net_15130), .Z(net_15131) );
SDFF_X2 inst_1347 ( .Q(net_8201), .D(net_8201), .SI(net_2713), .SE(net_2561), .CK(net_14431) );
SDFF_X2 inst_509 ( .Q(net_8862), .D(net_8862), .SI(net_3960), .SE(net_3936), .CK(net_13358) );
CLKBUF_X2 inst_11073 ( .A(net_10201), .Z(net_10921) );
SDFFR_X1 inst_2687 ( .SI(net_7549), .SE(net_5043), .CK(net_12753), .RN(x6501), .Q(x3938), .D(x3938) );
CLKBUF_X2 inst_11473 ( .A(net_11320), .Z(net_11321) );
CLKBUF_X2 inst_11775 ( .A(net_11241), .Z(net_11623) );
DFFR_X2 inst_7139 ( .QN(net_6401), .D(net_2934), .CK(net_15689), .RN(x6501) );
SDFFR_X2 inst_2622 ( .Q(net_7393), .D(net_7393), .SE(net_1136), .CK(net_15798), .RN(x6501), .SI(x4496) );
XNOR2_X2 inst_153 ( .ZN(net_2032), .B(net_1949), .A(net_1948) );
NAND2_X2 inst_4856 ( .ZN(net_1509), .A2(net_887), .A1(net_170) );
CLKBUF_X2 inst_9751 ( .A(net_9199), .Z(net_9599) );
SDFF_X2 inst_1459 ( .SI(net_7279), .Q(net_7136), .D(net_7136), .SE(net_6279), .CK(net_14632) );
NAND2_X2 inst_4094 ( .ZN(net_5441), .A1(net_5248), .A2(net_5017) );
CLKBUF_X2 inst_10483 ( .A(net_10330), .Z(net_10331) );
XNOR2_X2 inst_209 ( .B(net_1508), .ZN(net_1466), .A(net_1465) );
INV_X4 inst_6068 ( .ZN(net_2724), .A(net_159) );
SDFF_X2 inst_1781 ( .D(net_7287), .SI(net_6944), .Q(net_6944), .SE(net_6281), .CK(net_14896) );
INV_X2 inst_6365 ( .ZN(net_1892), .A(net_1891) );
CLKBUF_X2 inst_16304 ( .A(net_13560), .Z(net_16152) );
SDFFR_X1 inst_2769 ( .Q(net_7298), .SI(net_7262), .D(net_2127), .SE(net_1327), .CK(net_18246), .RN(x6501) );
CLKBUF_X2 inst_17794 ( .A(net_17641), .Z(net_17642) );
CLKBUF_X2 inst_17625 ( .A(net_17472), .Z(net_17473) );
INV_X2 inst_6230 ( .ZN(net_5480), .A(net_5306) );
CLKBUF_X2 inst_11353 ( .A(net_11200), .Z(net_11201) );
CLKBUF_X2 inst_15797 ( .A(net_15644), .Z(net_15645) );
NAND3_X2 inst_3982 ( .ZN(net_2004), .A3(net_1718), .A2(net_971), .A1(net_941) );
INV_X2 inst_6482 ( .A(net_5949), .ZN(net_895) );
OAI211_X2 inst_3215 ( .ZN(net_1746), .C1(net_1745), .B(net_1437), .A(net_1024), .C2(net_188) );
CLKBUF_X2 inst_14273 ( .A(net_12250), .Z(net_14121) );
CLKBUF_X2 inst_18231 ( .A(net_13338), .Z(net_18079) );
INV_X4 inst_5810 ( .A(net_7517), .ZN(net_1262) );
AOI22_X2 inst_8462 ( .B1(net_6653), .A1(net_6620), .A2(net_6213), .B2(net_6138), .ZN(net_3478) );
NAND2_X2 inst_4167 ( .ZN(net_5344), .A1(net_5089), .A2(net_5088) );
AND2_X2 inst_9204 ( .A1(net_7261), .ZN(net_898), .A2(net_897) );
NAND2_X2 inst_4374 ( .A1(net_7155), .A2(net_5166), .ZN(net_5083) );
SDFF_X2 inst_1995 ( .SI(net_7916), .Q(net_7916), .D(net_2702), .SE(net_2461), .CK(net_18029) );
CLKBUF_X2 inst_15031 ( .A(net_14878), .Z(net_14879) );
AND2_X4 inst_9145 ( .ZN(net_1296), .A2(net_211), .A1(net_167) );
CLKBUF_X2 inst_17894 ( .A(net_17741), .Z(net_17742) );
DFFR_X1 inst_7405 ( .D(net_5693), .CK(net_14047), .RN(x6501), .Q(x394) );
NOR2_X2 inst_3367 ( .ZN(net_5558), .A1(net_5360), .A2(net_5359) );
CLKBUF_X2 inst_12736 ( .A(net_12583), .Z(net_12584) );
SDFF_X2 inst_568 ( .Q(net_8832), .D(net_8832), .SI(net_3967), .SE(net_3964), .CK(net_13129) );
SDFF_X2 inst_523 ( .Q(net_8878), .D(net_8878), .SI(net_3975), .SE(net_3936), .CK(net_12543) );
SDFF_X2 inst_1483 ( .SI(net_7281), .Q(net_7098), .D(net_7098), .SE(net_6278), .CK(net_19030) );
CLKBUF_X2 inst_15445 ( .A(net_15292), .Z(net_15293) );
CLKBUF_X2 inst_17843 ( .A(net_12008), .Z(net_17691) );
CLKBUF_X2 inst_10202 ( .A(net_10049), .Z(net_10050) );
SDFF_X2 inst_1492 ( .SI(net_7293), .Q(net_7070), .D(net_7070), .SE(net_6280), .CK(net_18397) );
CLKBUF_X2 inst_18328 ( .A(net_13342), .Z(net_18176) );
NAND2_X2 inst_4234 ( .A1(net_7020), .A2(net_5249), .ZN(net_5226) );
DFF_X1 inst_6722 ( .Q(net_6768), .D(net_5647), .CK(net_9340) );
CLKBUF_X2 inst_11982 ( .A(net_11829), .Z(net_11830) );
CLKBUF_X2 inst_19061 ( .A(net_18908), .Z(net_18909) );
CLKBUF_X2 inst_16694 ( .A(net_16541), .Z(net_16542) );
OR2_X2 inst_2898 ( .A2(net_2739), .A1(net_599), .ZN(x4234) );
AOI21_X2 inst_8875 ( .ZN(net_5872), .B2(net_5871), .A(net_5844), .B1(x208) );
CLKBUF_X2 inst_10280 ( .A(net_10127), .Z(net_10128) );
CLKBUF_X2 inst_17162 ( .A(net_17009), .Z(net_17010) );
SDFF_X2 inst_1368 ( .SI(net_7280), .Q(net_7137), .D(net_7137), .SE(net_6279), .CK(net_19047) );
CLKBUF_X2 inst_13708 ( .A(net_13555), .Z(net_13556) );
CLKBUF_X2 inst_15665 ( .A(net_15512), .Z(net_15513) );
DFFR_X2 inst_7282 ( .QN(net_6389), .D(net_1774), .CK(net_15657), .RN(x6501) );
SDFFS_X2 inst_2088 ( .SI(net_6821), .Q(net_6821), .SE(net_2146), .D(net_1394), .CK(net_18684), .SN(x6501) );
DFF_X1 inst_6775 ( .Q(net_7554), .D(net_4597), .CK(net_12758) );
CLKBUF_X2 inst_15199 ( .A(net_15046), .Z(net_15047) );
CLKBUF_X2 inst_18565 ( .A(net_18412), .Z(net_18413) );
CLKBUF_X2 inst_17475 ( .A(net_15753), .Z(net_17323) );
CLKBUF_X2 inst_16026 ( .A(net_15873), .Z(net_15874) );
HA_X1 inst_6673 ( .S(net_3196), .CO(net_3195), .A(net_3194), .B(net_3015) );
SDFF_X2 inst_1379 ( .SI(net_7266), .Q(net_7123), .D(net_7123), .SE(net_6279), .CK(net_14375) );
CLKBUF_X2 inst_12326 ( .A(net_12173), .Z(net_12174) );
CLKBUF_X2 inst_9582 ( .A(net_9197), .Z(net_9430) );
CLKBUF_X2 inst_15739 ( .A(net_13170), .Z(net_15587) );
CLKBUF_X2 inst_12217 ( .A(net_12064), .Z(net_12065) );
CLKBUF_X2 inst_9221 ( .A(net_9068), .Z(net_9069) );
CLKBUF_X2 inst_15582 ( .A(net_15429), .Z(net_15430) );
INV_X4 inst_6131 ( .A(net_8925), .ZN(net_2610) );
CLKBUF_X2 inst_13643 ( .A(net_13490), .Z(net_13491) );
INV_X4 inst_5796 ( .A(net_7499), .ZN(net_3051) );
CLKBUF_X2 inst_14229 ( .A(net_14076), .Z(net_14077) );
CLKBUF_X2 inst_9571 ( .A(net_9418), .Z(net_9419) );
CLKBUF_X2 inst_14654 ( .A(net_12954), .Z(net_14502) );
CLKBUF_X2 inst_14924 ( .A(net_14771), .Z(net_14772) );
SDFF_X2 inst_583 ( .Q(net_8850), .D(net_8850), .SE(net_3964), .SI(net_3949), .CK(net_12618) );
SDFF_X2 inst_1904 ( .D(net_7266), .SI(net_7003), .Q(net_7003), .SE(net_6277), .CK(net_17055) );
CLKBUF_X2 inst_13970 ( .A(net_13817), .Z(net_13818) );
CLKBUF_X2 inst_10732 ( .A(net_10579), .Z(net_10580) );
CLKBUF_X2 inst_18156 ( .A(net_18003), .Z(net_18004) );
NAND2_X2 inst_4325 ( .A1(net_7041), .A2(net_5162), .ZN(net_5132) );
CLKBUF_X2 inst_10932 ( .A(net_9813), .Z(net_10780) );
CLKBUF_X2 inst_14146 ( .A(net_13993), .Z(net_13994) );
CLKBUF_X2 inst_10441 ( .A(net_10288), .Z(net_10289) );
DFFS_X1 inst_6913 ( .Q(net_6331), .D(net_5727), .CK(net_14213), .SN(x6501) );
DFF_X1 inst_6788 ( .Q(net_7644), .D(net_4591), .CK(net_10800) );
CLKBUF_X2 inst_17583 ( .A(net_9846), .Z(net_17431) );
CLKBUF_X2 inst_14346 ( .A(net_14193), .Z(net_14194) );
NAND2_X2 inst_4863 ( .A2(net_7346), .ZN(net_5986), .A1(net_844) );
NAND2_X1 inst_4910 ( .A1(net_8945), .ZN(net_1044), .A2(net_1043) );
CLKBUF_X2 inst_12513 ( .A(net_12360), .Z(net_12361) );
CLKBUF_X2 inst_14667 ( .A(net_14514), .Z(net_14515) );
CLKBUF_X2 inst_12113 ( .A(net_11960), .Z(net_11961) );
CLKBUF_X2 inst_14985 ( .A(net_14832), .Z(net_14833) );
CLKBUF_X2 inst_9811 ( .A(net_9658), .Z(net_9659) );
CLKBUF_X2 inst_14504 ( .A(net_14351), .Z(net_14352) );
CLKBUF_X2 inst_17523 ( .A(net_17370), .Z(net_17371) );
AOI222_X1 inst_8693 ( .C2(net_5832), .A2(net_5830), .B2(net_5824), .ZN(net_3210), .B1(net_2126), .A1(net_1775), .C1(x3418) );
INV_X4 inst_6025 ( .A(net_6354), .ZN(net_507) );
CLKBUF_X2 inst_17330 ( .A(net_17177), .Z(net_17178) );
SDFFR_X2 inst_2289 ( .SE(net_2436), .SI(net_2435), .Q(net_268), .D(net_268), .CK(net_16547), .RN(x6501) );
CLKBUF_X2 inst_18850 ( .A(net_18692), .Z(net_18698) );
SDFFR_X1 inst_2750 ( .SI(net_9029), .Q(net_9029), .D(net_7458), .SE(net_3208), .CK(net_10637), .RN(x6501) );
SDFF_X2 inst_1467 ( .SI(net_7265), .Q(net_7122), .D(net_7122), .SE(net_6279), .CK(net_17075) );
INV_X4 inst_5800 ( .A(net_7228), .ZN(net_1854) );
CLKBUF_X2 inst_14313 ( .A(net_14160), .Z(net_14161) );
INV_X4 inst_5772 ( .A(net_9010), .ZN(net_722) );
CLKBUF_X2 inst_10258 ( .A(net_10105), .Z(net_10106) );
CLKBUF_X2 inst_10803 ( .A(net_9208), .Z(net_10651) );
CLKBUF_X2 inst_14102 ( .A(net_13949), .Z(net_13950) );
INV_X2 inst_6317 ( .ZN(net_3346), .A(net_3291) );
CLKBUF_X2 inst_13227 ( .A(net_13074), .Z(net_13075) );
OR2_X4 inst_2834 ( .A1(net_6171), .ZN(net_3033), .A2(net_2849) );
CLKBUF_X2 inst_15067 ( .A(net_9109), .Z(net_14915) );
CLKBUF_X2 inst_17653 ( .A(net_17500), .Z(net_17501) );
CLKBUF_X2 inst_16064 ( .A(net_15911), .Z(net_15912) );
AOI22_X2 inst_8130 ( .B1(net_7913), .A1(net_7811), .B2(net_6103), .A2(net_4398), .ZN(net_4019) );
SDFF_X2 inst_1513 ( .SI(net_7844), .Q(net_7844), .D(net_2709), .SE(net_2558), .CK(net_15284) );
CLKBUF_X2 inst_9864 ( .A(net_9066), .Z(net_9712) );
CLKBUF_X2 inst_11756 ( .A(net_11603), .Z(net_11604) );
CLKBUF_X2 inst_10916 ( .A(net_10763), .Z(net_10764) );
NAND2_X2 inst_4080 ( .A2(net_6783), .A1(net_5835), .ZN(net_5766) );
CLKBUF_X2 inst_10846 ( .A(net_10693), .Z(net_10694) );
SDFF_X2 inst_1545 ( .Q(net_8001), .D(net_8001), .SI(net_2711), .SE(net_2542), .CK(net_17008) );
CLKBUF_X2 inst_12750 ( .A(net_12597), .Z(net_12598) );
NOR2_X4 inst_3338 ( .A1(net_7307), .ZN(net_1635), .A2(net_1524) );
SDFF_X2 inst_406 ( .SI(net_8319), .Q(net_8319), .SE(net_3978), .D(net_3963), .CK(net_12356) );
NAND2_X2 inst_4579 ( .A2(net_4362), .ZN(net_2958), .A1(net_2957) );
INV_X4 inst_5933 ( .A(net_7304), .ZN(net_655) );
CLKBUF_X2 inst_14696 ( .A(net_14543), .Z(net_14544) );
CLKBUF_X2 inst_13818 ( .A(net_13665), .Z(net_13666) );
XNOR2_X2 inst_328 ( .B(net_1026), .A(net_978), .ZN(net_924) );
CLKBUF_X2 inst_18677 ( .A(net_15465), .Z(net_18525) );
NAND2_X2 inst_4217 ( .A1(net_6892), .A2(net_5247), .ZN(net_5243) );
AOI22_X2 inst_8496 ( .B1(net_6547), .A1(net_6514), .A2(net_6137), .B2(net_6104), .ZN(net_3444) );
SDFF_X2 inst_818 ( .SI(net_8510), .Q(net_8510), .D(net_3953), .SE(net_3884), .CK(net_10231) );
CLKBUF_X2 inst_12373 ( .A(net_12220), .Z(net_12221) );
CLKBUF_X2 inst_18336 ( .A(net_18183), .Z(net_18184) );
CLKBUF_X2 inst_18229 ( .A(net_9157), .Z(net_18077) );
CLKBUF_X2 inst_9902 ( .A(net_9553), .Z(net_9750) );
CLKBUF_X2 inst_16959 ( .A(net_16806), .Z(net_16807) );
DFFR_X1 inst_7561 ( .D(net_7668), .Q(net_7656), .CK(net_12704), .RN(x6501) );
CLKBUF_X2 inst_9825 ( .A(net_9221), .Z(net_9673) );
CLKBUF_X2 inst_10172 ( .A(net_10019), .Z(net_10020) );
NOR3_X2 inst_3274 ( .A1(net_2415), .ZN(net_2412), .A3(net_2397), .A2(net_1090) );
CLKBUF_X2 inst_13920 ( .A(net_10453), .Z(net_13768) );
CLKBUF_X2 inst_11776 ( .A(net_11623), .Z(net_11624) );
CLKBUF_X2 inst_12643 ( .A(net_12490), .Z(net_12491) );
CLKBUF_X2 inst_17011 ( .A(net_16858), .Z(net_16859) );
AND2_X2 inst_9178 ( .ZN(net_2502), .A2(net_2241), .A1(net_574) );
CLKBUF_X2 inst_17207 ( .A(net_17054), .Z(net_17055) );
CLKBUF_X2 inst_10066 ( .A(net_9366), .Z(net_9914) );
AOI22_X2 inst_8360 ( .B1(net_8887), .A1(net_8332), .B2(net_6252), .A2(net_4345), .ZN(net_3688) );
CLKBUF_X2 inst_19151 ( .A(net_18998), .Z(net_18999) );
INV_X2 inst_6442 ( .ZN(net_618), .A(net_617) );
CLKBUF_X2 inst_15622 ( .A(net_10646), .Z(net_15470) );
CLKBUF_X2 inst_16850 ( .A(net_14129), .Z(net_16698) );
DFFR_X2 inst_7146 ( .QN(net_7365), .D(net_2886), .CK(net_11841), .RN(x6501) );
CLKBUF_X2 inst_16056 ( .A(net_15903), .Z(net_15904) );
SDFF_X2 inst_906 ( .SI(net_8705), .Q(net_8705), .SE(net_6195), .D(net_3943), .CK(net_13083) );
NAND2_X2 inst_4276 ( .A1(net_7003), .A2(net_5249), .ZN(net_5184) );
CLKBUF_X2 inst_17293 ( .A(net_12997), .Z(net_17141) );
INV_X4 inst_5222 ( .ZN(net_2678), .A(net_2220) );
INV_X4 inst_5098 ( .ZN(net_5695), .A(net_5667) );
CLKBUF_X2 inst_13600 ( .A(net_13447), .Z(net_13448) );
CLKBUF_X2 inst_16478 ( .A(net_16325), .Z(net_16326) );
SDFFR_X2 inst_2598 ( .QN(net_7246), .D(net_2803), .SI(net_1867), .SE(net_1379), .CK(net_18106), .RN(x6501) );
SDFF_X2 inst_1248 ( .SI(net_7692), .Q(net_7692), .SE(net_2714), .D(net_2712), .CK(net_17158) );
CLKBUF_X2 inst_18626 ( .A(net_18473), .Z(net_18474) );
NAND3_X2 inst_3998 ( .A3(net_2913), .A2(net_2827), .ZN(net_1497), .A1(net_1496) );
CLKBUF_X2 inst_18124 ( .A(net_12232), .Z(net_17972) );
CLKBUF_X2 inst_18867 ( .A(net_18714), .Z(net_18715) );
AND4_X2 inst_9035 ( .ZN(net_5284), .A4(net_4906), .A2(net_4582), .A3(net_4558), .A1(net_4496) );
CLKBUF_X2 inst_18779 ( .A(net_18626), .Z(net_18627) );
NAND2_X2 inst_4300 ( .A1(net_7092), .A2(net_5164), .ZN(net_5157) );
CLKBUF_X2 inst_12000 ( .A(net_10559), .Z(net_11848) );
CLKBUF_X2 inst_16221 ( .A(net_16068), .Z(net_16069) );
XNOR2_X2 inst_183 ( .ZN(net_1671), .B(net_1583), .A(net_1582) );
AOI22_X2 inst_7748 ( .B1(net_6977), .A1(net_6937), .A2(net_5443), .B2(net_5442), .ZN(net_5414) );
HA_X1 inst_6703 ( .CO(net_6188), .A(net_6176), .S(net_2149), .B(x3372) );
AOI22_X2 inst_8471 ( .B1(net_6607), .A1(net_6574), .A2(net_6257), .B2(net_6110), .ZN(net_3469) );
CLKBUF_X2 inst_15822 ( .A(net_12825), .Z(net_15670) );
CLKBUF_X2 inst_17266 ( .A(net_15117), .Z(net_17114) );
AOI22_X2 inst_8081 ( .B1(net_8046), .A1(net_7842), .B2(net_6107), .A2(net_4400), .ZN(net_4064) );
SDFF_X2 inst_1848 ( .D(net_7266), .SI(net_6883), .Q(net_6883), .SE(net_6284), .CK(net_14344) );
CLKBUF_X2 inst_12694 ( .A(net_12541), .Z(net_12542) );
NAND2_X2 inst_4451 ( .ZN(net_4975), .A2(net_4824), .A1(net_4485) );
SDFF_X2 inst_487 ( .SI(net_8611), .Q(net_8611), .SE(net_3984), .D(net_3958), .CK(net_10025) );
CLKBUF_X2 inst_11338 ( .A(net_11185), .Z(net_11186) );
CLKBUF_X2 inst_14540 ( .A(net_12818), .Z(net_14388) );
CLKBUF_X2 inst_17810 ( .A(net_17657), .Z(net_17658) );
INV_X4 inst_5315 ( .ZN(net_1681), .A(net_1129) );
CLKBUF_X2 inst_13696 ( .A(net_12351), .Z(net_13544) );
CLKBUF_X2 inst_17376 ( .A(net_17223), .Z(net_17224) );
SDFFR_X2 inst_2133 ( .SI(net_7201), .Q(net_7201), .D(net_6452), .SE(net_4362), .CK(net_13732), .RN(x6501) );
SDFFR_X2 inst_2163 ( .QN(net_7583), .D(net_3963), .SE(net_3144), .SI(net_3137), .CK(net_12656), .RN(x6501) );
CLKBUF_X2 inst_17882 ( .A(net_17729), .Z(net_17730) );
CLKBUF_X2 inst_19011 ( .A(net_9253), .Z(net_18859) );
CLKBUF_X2 inst_9947 ( .A(net_9794), .Z(net_9795) );
INV_X4 inst_6051 ( .A(net_8897), .ZN(net_496) );
NAND2_X2 inst_4668 ( .A2(net_6217), .A1(net_6216), .ZN(net_2239) );
INV_X4 inst_5497 ( .ZN(net_885), .A(net_713) );
SDFF_X2 inst_1861 ( .D(net_7292), .SI(net_6949), .Q(net_6949), .SE(net_6281), .CK(net_14882) );
NOR2_X2 inst_3570 ( .A2(net_6753), .ZN(net_2904), .A1(net_498) );
AND2_X4 inst_9133 ( .ZN(net_1389), .A2(net_814), .A1(net_175) );
NAND2_X2 inst_4835 ( .ZN(net_989), .A1(net_774), .A2(net_605) );
CLKBUF_X2 inst_15050 ( .A(net_14897), .Z(net_14898) );
OR2_X4 inst_2857 ( .A2(net_8950), .A1(net_8949), .ZN(net_619) );
AOI222_X1 inst_8667 ( .B1(net_7667), .A2(net_3599), .B2(net_3598), .C2(net_3597), .ZN(net_3591), .C1(net_1553), .A1(net_1358) );
CLKBUF_X2 inst_15116 ( .A(net_14963), .Z(net_14964) );
SDFF_X2 inst_1585 ( .Q(net_8039), .D(net_8039), .SI(net_2660), .SE(net_2545), .CK(net_16992) );
CLKBUF_X2 inst_10754 ( .A(net_10601), .Z(net_10602) );
CLKBUF_X2 inst_11412 ( .A(net_11259), .Z(net_11260) );
SDFF_X2 inst_1873 ( .D(net_7276), .SI(net_6973), .Q(net_6973), .SE(net_6283), .CK(net_17352) );
CLKBUF_X2 inst_11965 ( .A(net_11812), .Z(net_11813) );
AOI22_X2 inst_7854 ( .A2(net_5595), .B2(net_4881), .ZN(net_4653), .A1(net_325), .B1(net_243) );
INV_X4 inst_6135 ( .A(net_6295), .ZN(net_2736) );
CLKBUF_X2 inst_11765 ( .A(net_11612), .Z(net_11613) );
INV_X4 inst_5263 ( .A(net_2304), .ZN(net_2250) );
OAI21_X2 inst_3114 ( .B1(net_6420), .B2(net_2433), .ZN(net_2432), .A(net_2431) );
NOR2_X2 inst_3577 ( .A2(net_6413), .ZN(net_1102), .A1(net_564) );
CLKBUF_X2 inst_9451 ( .A(net_9298), .Z(net_9299) );
CLKBUF_X2 inst_15035 ( .A(net_9541), .Z(net_14883) );
NAND2_X2 inst_4754 ( .ZN(net_2717), .A1(net_1776), .A2(net_1586) );
CLKBUF_X2 inst_17711 ( .A(net_17558), .Z(net_17559) );
CLKBUF_X2 inst_10216 ( .A(net_9602), .Z(net_10064) );
CLKBUF_X2 inst_11554 ( .A(net_11401), .Z(net_11402) );
NAND2_X2 inst_4680 ( .ZN(net_2319), .A2(net_2082), .A1(net_2070) );
INV_X2 inst_6589 ( .A(net_6119), .ZN(net_6118) );
CLKBUF_X2 inst_16216 ( .A(net_16063), .Z(net_16064) );
CLKBUF_X2 inst_16952 ( .A(net_16799), .Z(net_16800) );
CLKBUF_X2 inst_14759 ( .A(net_14606), .Z(net_14607) );
SDFF_X2 inst_1727 ( .Q(net_7995), .D(net_7995), .SI(net_2722), .SE(net_2542), .CK(net_17690) );
SDFF_X2 inst_1753 ( .Q(net_8125), .D(net_8125), .SI(net_2720), .SE(net_2541), .CK(net_15233) );
SDFF_X2 inst_1166 ( .D(net_7314), .SI(net_6490), .Q(net_6490), .SE(net_3071), .CK(net_9896) );
XNOR2_X2 inst_116 ( .ZN(net_3201), .A(net_3047), .B(x2261) );
INV_X4 inst_5498 ( .A(net_1039), .ZN(net_709) );
INV_X2 inst_6559 ( .A(net_7567), .ZN(net_3131) );
CLKBUF_X2 inst_15183 ( .A(net_15030), .Z(net_15031) );
CLKBUF_X2 inst_10142 ( .A(net_9989), .Z(net_9990) );
NAND2_X2 inst_4087 ( .A1(net_6125), .ZN(net_5534), .A2(net_5533) );
SDFF_X2 inst_471 ( .SI(net_8476), .Q(net_8476), .SE(net_3983), .D(net_3951), .CK(net_10606) );
CLKBUF_X2 inst_10680 ( .A(net_10527), .Z(net_10528) );
CLKBUF_X2 inst_12104 ( .A(net_10246), .Z(net_11952) );
INV_X2 inst_6557 ( .A(net_7500), .ZN(net_497) );
CLKBUF_X2 inst_11081 ( .A(net_10130), .Z(net_10929) );
CLKBUF_X2 inst_18349 ( .A(net_18196), .Z(net_18197) );
SDFF_X2 inst_896 ( .SI(net_8713), .Q(net_8713), .SE(net_6195), .D(net_3946), .CK(net_10692) );
CLKBUF_X2 inst_12315 ( .A(net_12162), .Z(net_12163) );
CLKBUF_X2 inst_9276 ( .A(net_9123), .Z(net_9124) );
CLKBUF_X2 inst_14552 ( .A(net_14136), .Z(net_14400) );
CLKBUF_X2 inst_9317 ( .A(net_9164), .Z(net_9165) );
CLKBUF_X2 inst_15021 ( .A(net_14868), .Z(net_14869) );
DFFR_X1 inst_7445 ( .QN(net_8925), .D(net_4758), .CK(net_13968), .RN(x6501) );
AOI22_X2 inst_8577 ( .B1(net_2571), .ZN(net_1590), .A1(net_1589), .A2(net_1588), .B2(net_1517) );
SDFFR_X2 inst_2557 ( .QN(net_6355), .SE(net_2147), .SI(net_1856), .D(net_727), .CK(net_17531), .RN(x6501) );
DFFR_X1 inst_7438 ( .QN(net_8936), .D(net_4746), .CK(net_14595), .RN(x6501) );
CLKBUF_X2 inst_15639 ( .A(net_13415), .Z(net_15487) );
NOR3_X2 inst_3319 ( .ZN(net_4469), .A3(net_1633), .A1(net_1431), .A2(net_1267) );
CLKBUF_X2 inst_15718 ( .A(net_15565), .Z(net_15566) );
NAND2_X2 inst_4621 ( .A2(net_6144), .ZN(net_2599), .A1(net_2598) );
CLKBUF_X2 inst_11519 ( .A(net_11366), .Z(net_11367) );
CLKBUF_X2 inst_17262 ( .A(net_13929), .Z(net_17110) );
SDFFR_X2 inst_2550 ( .QN(net_6367), .SE(net_2147), .D(net_2134), .SI(net_1955), .CK(net_14748), .RN(x6501) );
CLKBUF_X2 inst_18826 ( .A(net_10712), .Z(net_18674) );
CLKBUF_X2 inst_14966 ( .A(net_14813), .Z(net_14814) );
CLKBUF_X2 inst_16301 ( .A(net_16148), .Z(net_16149) );
DFFR_X1 inst_7559 ( .D(net_6483), .Q(net_6465), .CK(net_15129), .RN(x6501) );
NAND2_X2 inst_4281 ( .A1(net_6885), .A2(net_5247), .ZN(net_5179) );
SDFFR_X2 inst_2142 ( .SI(net_7181), .Q(net_7181), .D(net_6432), .SE(net_4362), .CK(net_13553), .RN(x6501) );
CLKBUF_X2 inst_16425 ( .A(net_9178), .Z(net_16273) );
CLKBUF_X2 inst_12810 ( .A(net_12657), .Z(net_12658) );
CLKBUF_X2 inst_18021 ( .A(net_17868), .Z(net_17869) );
INV_X4 inst_5110 ( .ZN(net_4946), .A(net_4879) );
DFF_X1 inst_6817 ( .QN(net_8229), .D(net_4452), .CK(net_17213) );
CLKBUF_X2 inst_19021 ( .A(net_18868), .Z(net_18869) );
NAND2_X2 inst_4458 ( .ZN(net_4934), .A2(net_4713), .A1(net_4495) );
CLKBUF_X2 inst_9407 ( .A(net_9058), .Z(net_9255) );
CLKBUF_X2 inst_14055 ( .A(net_11191), .Z(net_13903) );
INV_X4 inst_5184 ( .A(net_4850), .ZN(net_4764) );
CLKBUF_X2 inst_10518 ( .A(net_10365), .Z(net_10366) );
CLKBUF_X2 inst_15767 ( .A(net_15614), .Z(net_15615) );
SDFF_X2 inst_547 ( .Q(net_8691), .D(net_8691), .SI(net_3955), .SE(net_3935), .CK(net_11015) );
AND2_X4 inst_9107 ( .ZN(net_2038), .A2(net_2037), .A1(net_523) );
CLKBUF_X2 inst_16399 ( .A(net_12861), .Z(net_16247) );
SDFF_X2 inst_1607 ( .Q(net_8143), .D(net_8143), .SI(net_2716), .SE(net_2541), .CK(net_16824) );
CLKBUF_X2 inst_11847 ( .A(net_11694), .Z(net_11695) );
CLKBUF_X2 inst_10367 ( .A(net_10214), .Z(net_10215) );
CLKBUF_X2 inst_11623 ( .A(net_9278), .Z(net_11471) );
SDFF_X2 inst_1854 ( .D(net_7280), .SI(net_6937), .Q(net_6937), .SE(net_6281), .CK(net_18991) );
AOI21_X2 inst_9002 ( .B1(net_6324), .B2(net_2309), .ZN(net_2179), .A(net_1061) );
CLKBUF_X2 inst_12676 ( .A(net_12523), .Z(net_12524) );
SDFF_X2 inst_1710 ( .Q(net_8121), .D(net_8121), .SI(net_2573), .SE(net_2541), .CK(net_15251) );
INV_X4 inst_5922 ( .A(net_6362), .ZN(net_525) );
DFFR_X2 inst_7295 ( .Q(net_7623), .D(net_1181), .CK(net_11142), .RN(x6501) );
CLKBUF_X2 inst_18748 ( .A(net_15160), .Z(net_18596) );
SDFFR_X2 inst_2407 ( .SE(net_2260), .Q(net_319), .D(net_319), .CK(net_10403), .RN(x6501), .SI(x3156) );
NAND2_X2 inst_4884 ( .A2(net_7348), .A1(net_7347), .ZN(net_1063) );
CLKBUF_X2 inst_13814 ( .A(net_12626), .Z(net_13662) );
OAI21_X2 inst_3142 ( .B2(net_2060), .ZN(net_2053), .A(net_1988), .B1(net_1347) );
DFFR_X1 inst_7516 ( .Q(net_6340), .D(net_1602), .CK(net_18969), .RN(x6501) );
SDFF_X2 inst_753 ( .Q(net_8793), .D(net_8793), .SI(net_3973), .SE(net_3879), .CK(net_12335) );
CLKBUF_X2 inst_9647 ( .A(net_9456), .Z(net_9495) );
NOR2_X2 inst_3427 ( .A2(net_3093), .ZN(net_3085), .A1(net_2036) );
INV_X4 inst_5486 ( .ZN(net_2277), .A(net_731) );
INV_X2 inst_6262 ( .A(net_8241), .ZN(net_4635) );
INV_X4 inst_5768 ( .A(net_7514), .ZN(net_661) );
DFFS_X1 inst_6946 ( .D(net_6145), .CK(net_16343), .SN(x6501), .Q(x886) );
SDFF_X2 inst_1954 ( .D(net_7263), .SI(net_7000), .Q(net_7000), .SE(net_6277), .CK(net_17049) );
NAND3_X2 inst_3941 ( .ZN(net_4836), .A2(net_4554), .A3(net_4553), .A1(net_1814) );
CLKBUF_X2 inst_16484 ( .A(net_16221), .Z(net_16332) );
AOI22_X2 inst_7815 ( .A2(net_8221), .B2(net_6144), .A1(net_4764), .ZN(net_4739), .B1(net_4669) );
CLKBUF_X2 inst_13543 ( .A(net_13390), .Z(net_13391) );
CLKBUF_X2 inst_10588 ( .A(net_10435), .Z(net_10436) );
CLKBUF_X2 inst_12746 ( .A(net_12003), .Z(net_12594) );
NAND4_X2 inst_3858 ( .A2(net_3990), .A1(net_3581), .ZN(net_1440), .A3(net_591), .A4(net_528) );
DFFR_X2 inst_7014 ( .QN(net_6310), .D(net_5744), .CK(net_16741), .RN(x6501) );
CLKBUF_X2 inst_13129 ( .A(net_12976), .Z(net_12977) );
CLKBUF_X2 inst_13949 ( .A(net_13796), .Z(net_13797) );
CLKBUF_X2 inst_13008 ( .A(net_10977), .Z(net_12856) );
DFFR_X2 inst_7342 ( .Q(net_7338), .CK(net_11716), .D(x12929), .RN(x6501) );
INV_X4 inst_5105 ( .ZN(net_5670), .A(net_5601) );
AOI221_X2 inst_8818 ( .B2(net_6441), .B1(net_5654), .A(net_4898), .C2(net_4881), .ZN(net_4681), .C1(net_241) );
CLKBUF_X2 inst_19057 ( .A(net_18904), .Z(net_18905) );
CLKBUF_X2 inst_18990 ( .A(net_16169), .Z(net_18838) );
CLKBUF_X2 inst_12725 ( .A(net_9680), .Z(net_12573) );
NOR2_X2 inst_3561 ( .A1(net_1657), .ZN(net_1326), .A2(net_1325) );
DFFR_X2 inst_7233 ( .QN(net_7360), .D(net_2194), .CK(net_11818), .RN(x6501) );
CLKBUF_X2 inst_17773 ( .A(net_9071), .Z(net_17621) );
CLKBUF_X2 inst_14286 ( .A(net_11237), .Z(net_14134) );
CLKBUF_X2 inst_18009 ( .A(net_17856), .Z(net_17857) );
OAI21_X2 inst_3046 ( .B2(net_8220), .B1(net_4928), .ZN(net_4773), .A(net_2937) );
AOI221_X2 inst_8751 ( .C2(net_6449), .C1(net_5654), .ZN(net_5596), .B2(net_5595), .A(net_5335), .B1(net_331) );
CLKBUF_X2 inst_16511 ( .A(net_16358), .Z(net_16359) );
NAND2_X2 inst_4644 ( .ZN(net_2443), .A2(net_2158), .A1(net_1769) );
NAND2_X2 inst_4844 ( .A1(net_7481), .A2(net_3921), .ZN(net_1325) );
CLKBUF_X2 inst_14994 ( .A(net_14841), .Z(net_14842) );
NAND4_X2 inst_3757 ( .ZN(net_4264), .A1(net_3848), .A2(net_3847), .A3(net_3846), .A4(net_3845) );
SDFF_X2 inst_917 ( .SI(net_8737), .Q(net_8737), .SE(net_6195), .D(net_3976), .CK(net_10310) );
NAND4_X2 inst_3712 ( .ZN(net_4425), .A4(net_4332), .A1(net_3687), .A2(net_3686), .A3(net_3685) );
SDFF_X2 inst_1743 ( .Q(net_7876), .D(net_7876), .SI(net_2705), .SE(net_2543), .CK(net_15815) );
CLKBUF_X2 inst_11713 ( .A(net_11560), .Z(net_11561) );
CLKBUF_X2 inst_13403 ( .A(net_13250), .Z(net_13251) );
XNOR2_X2 inst_215 ( .B(net_7166), .ZN(net_1428), .A(net_1427) );
INV_X8 inst_5022 ( .ZN(net_3936), .A(net_3364) );
SDFFR_X2 inst_2624 ( .Q(net_7387), .D(net_7387), .SE(net_1136), .CK(net_18302), .RN(x6501), .SI(x4576) );
CLKBUF_X2 inst_18524 ( .A(net_18371), .Z(net_18372) );
INV_X2 inst_6258 ( .ZN(net_4658), .A(net_4569) );
DFFR_X1 inst_7550 ( .Q(net_8265), .D(net_976), .CK(net_15704), .RN(x6501) );
CLKBUF_X2 inst_11293 ( .A(net_10536), .Z(net_11141) );
CLKBUF_X2 inst_17089 ( .A(net_16936), .Z(net_16937) );
CLKBUF_X2 inst_17060 ( .A(net_16907), .Z(net_16908) );
CLKBUF_X2 inst_15848 ( .A(net_13670), .Z(net_15696) );
AOI21_X2 inst_8912 ( .ZN(net_5807), .A(net_5745), .B2(net_5608), .B1(net_5257) );
CLKBUF_X2 inst_17901 ( .A(net_17748), .Z(net_17749) );
NAND2_X2 inst_4819 ( .A1(net_6322), .ZN(net_1374), .A2(net_860) );
CLKBUF_X2 inst_15437 ( .A(net_11329), .Z(net_15285) );
CLKBUF_X2 inst_17544 ( .A(net_17391), .Z(net_17392) );
CLKBUF_X2 inst_16927 ( .A(net_16774), .Z(net_16775) );
NAND2_X2 inst_4774 ( .A2(net_2528), .ZN(net_1711), .A1(net_1634) );
CLKBUF_X2 inst_12997 ( .A(net_12844), .Z(net_12845) );
AOI222_X1 inst_8622 ( .A2(net_8226), .A1(net_4891), .B2(net_4889), .C2(net_4888), .ZN(net_4883), .B1(net_4714), .C1(net_3130) );
CLKBUF_X2 inst_18060 ( .A(net_17907), .Z(net_17908) );
CLKBUF_X2 inst_12401 ( .A(net_12248), .Z(net_12249) );
CLKBUF_X2 inst_17454 ( .A(net_17301), .Z(net_17302) );
CLKBUF_X2 inst_18300 ( .A(net_12093), .Z(net_18148) );
CLKBUF_X2 inst_14632 ( .A(net_13119), .Z(net_14480) );
CLKBUF_X2 inst_18876 ( .A(net_9541), .Z(net_18724) );
NAND2_X4 inst_4016 ( .ZN(net_4415), .A1(net_4376), .A2(net_4356) );
OAI22_X2 inst_2914 ( .ZN(net_3970), .A2(net_3552), .B2(net_3549), .A1(net_1370), .B1(net_694) );
NOR3_X2 inst_3294 ( .ZN(net_2024), .A1(net_1834), .A3(net_1390), .A2(net_1388) );
SDFFR_X1 inst_2741 ( .SI(net_9024), .Q(net_9024), .D(net_7453), .SE(net_3208), .CK(net_12841), .RN(x6501) );
CLKBUF_X2 inst_11825 ( .A(net_11672), .Z(net_11673) );
CLKBUF_X2 inst_15262 ( .A(net_15109), .Z(net_15110) );
CLKBUF_X2 inst_11966 ( .A(net_11813), .Z(net_11814) );
SDFF_X2 inst_1522 ( .Q(net_7893), .D(net_7893), .SI(net_2722), .SE(net_2543), .CK(net_17698) );
CLKBUF_X2 inst_14380 ( .A(net_14227), .Z(net_14228) );
CLKBUF_X2 inst_12135 ( .A(net_11982), .Z(net_11983) );
CLKBUF_X2 inst_11455 ( .A(net_11302), .Z(net_11303) );
CLKBUF_X2 inst_13955 ( .A(net_13218), .Z(net_13803) );
CLKBUF_X2 inst_16931 ( .A(net_16778), .Z(net_16779) );
CLKBUF_X2 inst_18964 ( .A(net_18811), .Z(net_18812) );
AOI222_X1 inst_8645 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3923), .B1(net_3391), .C1(net_3390), .A1(x13698) );
CLKBUF_X2 inst_16566 ( .A(net_16413), .Z(net_16414) );
INV_X4 inst_5761 ( .A(net_5965), .ZN(x3079) );
DFFS_X1 inst_6964 ( .Q(net_8264), .D(net_956), .CK(net_18484), .SN(x6501) );
CLKBUF_X2 inst_12520 ( .A(net_10238), .Z(net_12368) );
CLKBUF_X2 inst_12809 ( .A(net_11649), .Z(net_12657) );
CLKBUF_X2 inst_9528 ( .A(net_9375), .Z(net_9376) );
CLKBUF_X2 inst_11889 ( .A(net_11736), .Z(net_11737) );
INV_X4 inst_5691 ( .ZN(net_2698), .A(net_143) );
AOI22_X2 inst_7902 ( .A2(net_5538), .ZN(net_4525), .B2(net_4388), .B1(net_2608), .A1(net_418) );
SDFF_X2 inst_861 ( .Q(net_8569), .D(net_8569), .SI(net_3966), .SE(net_3878), .CK(net_9980) );
AOI22_X2 inst_8392 ( .B1(net_8710), .A1(net_8488), .ZN(net_6071), .B2(net_4350), .A2(net_4349) );
CLKBUF_X2 inst_18937 ( .A(net_18784), .Z(net_18785) );
DFFR_X1 inst_7431 ( .QN(net_8938), .D(net_4856), .CK(net_16442), .RN(x6501) );
CLKBUF_X2 inst_11549 ( .A(net_11396), .Z(net_11397) );
OAI21_X2 inst_2990 ( .B2(net_5912), .ZN(net_5904), .A(net_5799), .B1(net_637) );
DFFR_X1 inst_7495 ( .QN(net_6399), .D(net_3092), .CK(net_15722), .RN(x6501) );
SDFF_X2 inst_1283 ( .Q(net_7832), .D(net_7832), .SE(net_2730), .SI(net_2710), .CK(net_16517) );
CLKBUF_X2 inst_17345 ( .A(net_9420), .Z(net_17193) );
CLKBUF_X2 inst_18299 ( .A(net_18146), .Z(net_18147) );
CLKBUF_X2 inst_11225 ( .A(net_11072), .Z(net_11073) );
CLKBUF_X2 inst_17232 ( .A(net_10258), .Z(net_17080) );
CLKBUF_X2 inst_10625 ( .A(net_10472), .Z(net_10473) );
NAND2_X2 inst_4290 ( .A1(net_7120), .ZN(net_5170), .A2(net_5166) );
CLKBUF_X2 inst_18050 ( .A(net_17897), .Z(net_17898) );
CLKBUF_X2 inst_16796 ( .A(net_16643), .Z(net_16644) );
CLKBUF_X2 inst_12594 ( .A(net_12441), .Z(net_12442) );
CLKBUF_X2 inst_11027 ( .A(net_10874), .Z(net_10875) );
CLKBUF_X2 inst_15104 ( .A(net_14951), .Z(net_14952) );
CLKBUF_X2 inst_17918 ( .A(net_17765), .Z(net_17766) );
CLKBUF_X2 inst_10238 ( .A(net_9280), .Z(net_10086) );
CLKBUF_X2 inst_16321 ( .A(net_16168), .Z(net_16169) );
INV_X4 inst_5195 ( .ZN(net_2861), .A(net_2664) );
CLKBUF_X2 inst_14701 ( .A(net_14548), .Z(net_14549) );
CLKBUF_X2 inst_18002 ( .A(net_17849), .Z(net_17850) );
CLKBUF_X2 inst_19044 ( .A(net_18891), .Z(net_18892) );
NOR2_X2 inst_3462 ( .A2(net_6135), .ZN(net_2804), .A1(net_1435) );
CLKBUF_X2 inst_16353 ( .A(net_16200), .Z(net_16201) );
NAND2_X2 inst_4254 ( .A1(net_7002), .A2(net_5249), .ZN(net_5206) );
AOI22_X2 inst_8288 ( .B1(net_8767), .A1(net_8397), .A2(net_3867), .B2(net_3866), .ZN(net_3754) );
NAND2_X2 inst_4330 ( .A1(net_7101), .A2(net_5164), .ZN(net_5127) );
CLKBUF_X2 inst_10031 ( .A(net_9878), .Z(net_9879) );
CLKBUF_X2 inst_11925 ( .A(net_11324), .Z(net_11773) );
CLKBUF_X2 inst_14220 ( .A(net_14067), .Z(net_14068) );
CLKBUF_X2 inst_19085 ( .A(net_10738), .Z(net_18933) );
CLKBUF_X2 inst_12204 ( .A(net_10527), .Z(net_12052) );
CLKBUF_X2 inst_9388 ( .A(net_9235), .Z(net_9236) );
SDFFR_X1 inst_2754 ( .QN(net_7574), .D(net_3966), .SE(net_3144), .SI(net_3142), .CK(net_13225), .RN(x6501) );
SDFF_X2 inst_794 ( .SI(net_8365), .Q(net_8365), .D(net_3951), .SE(net_3880), .CK(net_13397) );
CLKBUF_X2 inst_14577 ( .A(net_14424), .Z(net_14425) );
CLKBUF_X2 inst_17864 ( .A(net_17711), .Z(net_17712) );
DFFR_X2 inst_7354 ( .Q(net_7324), .CK(net_11765), .D(x13058), .RN(x6501) );
CLKBUF_X2 inst_17663 ( .A(net_17510), .Z(net_17511) );
CLKBUF_X2 inst_12049 ( .A(net_9968), .Z(net_11897) );
SDFFR_X1 inst_2759 ( .QN(net_7566), .D(net_3965), .SE(net_3144), .SI(net_3132), .CK(net_10796), .RN(x6501) );
CLKBUF_X2 inst_17378 ( .A(net_11306), .Z(net_17226) );
CLKBUF_X2 inst_12092 ( .A(net_11939), .Z(net_11940) );
AOI22_X2 inst_8256 ( .B1(net_8726), .A1(net_8504), .B2(net_4350), .A2(net_4349), .ZN(net_3782) );
CLKBUF_X2 inst_11165 ( .A(net_11012), .Z(net_11013) );
SDFFR_X2 inst_2423 ( .D(net_2679), .SE(net_2678), .SI(net_472), .Q(net_472), .CK(net_16906), .RN(x6501) );
CLKBUF_X2 inst_16131 ( .A(net_15978), .Z(net_15979) );
SDFF_X2 inst_996 ( .D(net_7335), .SI(net_6643), .Q(net_6643), .SE(net_3123), .CK(net_9765) );
CLKBUF_X2 inst_10963 ( .A(net_10810), .Z(net_10811) );
INV_X4 inst_5889 ( .A(net_7411), .ZN(net_2021) );
CLKBUF_X2 inst_16230 ( .A(net_16077), .Z(net_16078) );
CLKBUF_X2 inst_12074 ( .A(net_11095), .Z(net_11922) );
SDFF_X2 inst_1527 ( .Q(net_7902), .D(net_7902), .SI(net_2715), .SE(net_2543), .CK(net_14182) );
INV_X4 inst_6142 ( .A(net_6132), .ZN(net_6130) );
SDFF_X2 inst_740 ( .Q(net_8786), .D(net_8786), .SI(net_3937), .SE(net_3879), .CK(net_11058) );
NAND2_X2 inst_4189 ( .ZN(net_5312), .A2(net_5184), .A1(net_5066) );
AOI22_X2 inst_7803 ( .A2(net_8247), .A1(net_5268), .ZN(net_4771), .B1(net_4743), .B2(net_4388) );
CLKBUF_X2 inst_17324 ( .A(net_17024), .Z(net_17172) );
DFF_X1 inst_6803 ( .QN(net_8249), .D(net_4430), .CK(net_16267) );
SDFF_X2 inst_1937 ( .SI(net_8069), .Q(net_8069), .D(net_2711), .SE(net_2508), .CK(net_14245) );
CLKBUF_X2 inst_15756 ( .A(net_10085), .Z(net_15604) );
SDFF_X2 inst_611 ( .SI(net_8407), .Q(net_8407), .SE(net_3969), .D(net_3948), .CK(net_13411) );
NAND2_X2 inst_4405 ( .A1(net_7088), .A2(net_5164), .ZN(net_5052) );
CLKBUF_X2 inst_10550 ( .A(net_10397), .Z(net_10398) );
SDFFR_X2 inst_2487 ( .D(net_7367), .SE(net_2548), .SI(net_2547), .QN(net_260), .CK(net_13544), .RN(x6501) );
CLKBUF_X2 inst_12417 ( .A(net_10735), .Z(net_12265) );
CLKBUF_X2 inst_12462 ( .A(net_12309), .Z(net_12310) );
CLKBUF_X2 inst_12549 ( .A(net_12396), .Z(net_12397) );
CLKBUF_X2 inst_16622 ( .A(net_16469), .Z(net_16470) );
AOI22_X2 inst_7802 ( .A2(net_4965), .ZN(net_4777), .B2(net_4397), .B1(net_2001), .A1(net_388) );
CLKBUF_X2 inst_15856 ( .A(net_15703), .Z(net_15704) );
SDFF_X2 inst_490 ( .SI(net_8614), .Q(net_8614), .SE(net_3984), .D(net_3956), .CK(net_13273) );
DFFR_X2 inst_7305 ( .D(net_6480), .QN(net_6477), .CK(net_11724), .RN(x6501) );
AOI22_X2 inst_8375 ( .B1(net_8708), .A1(net_8486), .B2(net_4350), .A2(net_4349), .ZN(net_3673) );
CLKBUF_X2 inst_13378 ( .A(net_12507), .Z(net_13226) );
SDFFR_X2 inst_2218 ( .Q(net_7451), .D(net_7451), .SE(net_2863), .CK(net_12926), .SI(x13567), .RN(x6501) );
SDFF_X2 inst_1309 ( .SI(net_7679), .Q(net_7679), .SE(net_2714), .D(net_2573), .CK(net_15294) );
CLKBUF_X2 inst_18396 ( .A(net_10250), .Z(net_18244) );
CLKBUF_X2 inst_15045 ( .A(net_14892), .Z(net_14893) );
NAND4_X2 inst_3803 ( .ZN(net_3623), .A1(net_3475), .A2(net_3474), .A3(net_3473), .A4(net_3472) );
MUX2_X2 inst_4938 ( .S(net_2852), .Z(net_2851), .B(net_2430), .A(net_904) );
CLKBUF_X2 inst_15049 ( .A(net_9188), .Z(net_14897) );
CLKBUF_X2 inst_16103 ( .A(net_11929), .Z(net_15951) );
OAI211_X2 inst_3183 ( .C2(net_6132), .ZN(net_5285), .B(net_4882), .A(net_4571), .C1(net_1419) );
CLKBUF_X2 inst_10242 ( .A(net_10089), .Z(net_10090) );
CLKBUF_X2 inst_13234 ( .A(net_13081), .Z(net_13082) );
CLKBUF_X2 inst_15095 ( .A(net_14942), .Z(net_14943) );
CLKBUF_X2 inst_10860 ( .A(net_10707), .Z(net_10708) );
CLKBUF_X2 inst_16498 ( .A(net_16345), .Z(net_16346) );
CLKBUF_X2 inst_19079 ( .A(net_18926), .Z(net_18927) );
CLKBUF_X2 inst_13301 ( .A(net_13148), .Z(net_13149) );
NAND2_X2 inst_4312 ( .A1(net_7096), .A2(net_5164), .ZN(net_5145) );
CLKBUF_X2 inst_11256 ( .A(net_11103), .Z(net_11104) );
CLKBUF_X2 inst_12950 ( .A(net_12797), .Z(net_12798) );
INV_X4 inst_5328 ( .ZN(net_1813), .A(net_1479) );
AOI22_X2 inst_8410 ( .B1(net_8713), .A1(net_8491), .B2(net_4350), .A2(net_4349), .ZN(net_3642) );
INV_X2 inst_6226 ( .ZN(net_5484), .A(net_5322) );
CLKBUF_X2 inst_13161 ( .A(net_13008), .Z(net_13009) );
CLKBUF_X2 inst_18782 ( .A(net_18629), .Z(net_18630) );
XNOR2_X2 inst_300 ( .ZN(net_981), .A(net_980), .B(net_520) );
CLKBUF_X2 inst_15407 ( .A(net_15254), .Z(net_15255) );
SDFF_X2 inst_1226 ( .Q(net_7960), .D(net_7960), .SE(net_2755), .SI(net_2590), .CK(net_16012) );
INV_X4 inst_5964 ( .A(net_7566), .ZN(net_517) );
CLKBUF_X2 inst_17836 ( .A(net_12442), .Z(net_17684) );
SDFF_X2 inst_446 ( .Q(net_8776), .D(net_8776), .SE(net_3982), .SI(net_3949), .CK(net_12634) );
AOI221_X2 inst_8802 ( .B1(net_7190), .C2(net_6129), .B2(net_5655), .A(net_4905), .ZN(net_4832), .C1(net_1401) );
CLKBUF_X2 inst_15619 ( .A(net_15466), .Z(net_15467) );
CLKBUF_X2 inst_15949 ( .A(net_15796), .Z(net_15797) );
MUX2_X2 inst_4923 ( .S(net_6328), .Z(net_4489), .A(net_489), .B(x4295) );
CLKBUF_X2 inst_18689 ( .A(net_18536), .Z(net_18537) );
NOR2_X2 inst_3533 ( .ZN(net_2181), .A1(net_1129), .A2(net_716) );
SDFF_X2 inst_824 ( .SI(net_8517), .Q(net_8517), .D(net_3949), .SE(net_3884), .CK(net_12579) );
CLKBUF_X2 inst_15996 ( .A(net_9916), .Z(net_15844) );
AOI22_X2 inst_7839 ( .B2(net_5595), .A2(net_5267), .ZN(net_4672), .A1(net_4671), .B1(net_338) );
CLKBUF_X2 inst_12897 ( .A(net_9174), .Z(net_12745) );
CLKBUF_X2 inst_10393 ( .A(net_9883), .Z(net_10241) );
CLKBUF_X2 inst_14678 ( .A(net_14525), .Z(net_14526) );
CLKBUF_X2 inst_16135 ( .A(net_15982), .Z(net_15983) );
INV_X2 inst_6600 ( .A(net_6155), .ZN(net_6152) );
AOI211_X2 inst_9007 ( .C2(net_5655), .ZN(net_5459), .A(net_4951), .B(net_4829), .C1(net_2953) );
CLKBUF_X2 inst_13691 ( .A(net_13538), .Z(net_13539) );
NAND4_X2 inst_3750 ( .ZN(net_4280), .A1(net_4014), .A2(net_4013), .A3(net_4012), .A4(net_4011) );
CLKBUF_X2 inst_11173 ( .A(net_11020), .Z(net_11021) );
CLKBUF_X2 inst_15286 ( .A(net_15133), .Z(net_15134) );
NAND2_X2 inst_4056 ( .ZN(net_5928), .A2(net_5927), .A1(net_2513) );
NAND2_X2 inst_4401 ( .A1(net_7127), .A2(net_5166), .ZN(net_5056) );
NOR2_X2 inst_3430 ( .A2(net_6143), .ZN(net_3185), .A1(net_3080) );
CLKBUF_X2 inst_10388 ( .A(net_10235), .Z(net_10236) );
CLKBUF_X2 inst_13368 ( .A(net_13215), .Z(net_13216) );
INV_X4 inst_5462 ( .ZN(net_1253), .A(net_1252) );
NOR2_X2 inst_3439 ( .A2(net_3093), .ZN(net_3058), .A1(net_2878) );
CLKBUF_X2 inst_17159 ( .A(net_17006), .Z(net_17007) );
CLKBUF_X2 inst_13968 ( .A(net_13815), .Z(net_13816) );
INV_X4 inst_5412 ( .ZN(net_1136), .A(net_868) );
AOI22_X2 inst_8308 ( .B1(net_8807), .A1(net_8548), .A2(net_3861), .B2(net_3860), .ZN(net_3737) );
CLKBUF_X2 inst_10901 ( .A(net_10639), .Z(net_10749) );
CLKBUF_X2 inst_10014 ( .A(net_9861), .Z(net_9862) );
CLKBUF_X2 inst_12459 ( .A(net_12306), .Z(net_12307) );
INV_X2 inst_6601 ( .A(net_6157), .ZN(net_6156) );
AOI22_X2 inst_8520 ( .B1(net_6552), .A1(net_6519), .A2(net_6137), .B2(net_6104), .ZN(net_3420) );
SDFF_X2 inst_1571 ( .SI(net_7736), .Q(net_7736), .D(net_2656), .SE(net_2559), .CK(net_17140) );
CLKBUF_X2 inst_15540 ( .A(net_9723), .Z(net_15388) );
CLKBUF_X2 inst_12009 ( .A(net_10091), .Z(net_11857) );
CLKBUF_X2 inst_17446 ( .A(net_13755), .Z(net_17294) );
AOI22_X2 inst_8214 ( .B1(net_8683), .A1(net_8646), .B2(net_6109), .A2(net_3857), .ZN(net_3822) );
SDFF_X2 inst_1402 ( .Q(net_8210), .D(net_8210), .SI(net_2704), .SE(net_2561), .CK(net_14288) );
INV_X2 inst_6511 ( .A(net_7219), .ZN(net_1872) );
CLKBUF_X2 inst_11246 ( .A(net_10128), .Z(net_11094) );
OAI21_X2 inst_3106 ( .ZN(net_2492), .B2(net_2489), .A(net_2332), .B1(net_2040) );
DFF_X1 inst_6810 ( .QN(net_8227), .D(net_4418), .CK(net_16552) );
CLKBUF_X2 inst_18586 ( .A(net_18433), .Z(net_18434) );
DFF_X1 inst_6843 ( .Q(net_6433), .D(net_3604), .CK(net_17967) );
CLKBUF_X2 inst_13379 ( .A(net_13226), .Z(net_13227) );
CLKBUF_X2 inst_17366 ( .A(net_11976), .Z(net_17214) );
INV_X2 inst_6270 ( .A(net_8235), .ZN(net_4626) );
INV_X4 inst_5453 ( .A(net_3299), .ZN(net_796) );
INV_X4 inst_5405 ( .ZN(net_3546), .A(net_877) );
AOI221_X2 inst_8810 ( .B1(net_9003), .C2(net_5535), .B2(net_5456), .A(net_4898), .ZN(net_4718), .C1(net_475) );
CLKBUF_X2 inst_13317 ( .A(net_13164), .Z(net_13165) );
SDFFR_X2 inst_2503 ( .Q(net_8977), .D(net_8977), .SI(net_4666), .SE(net_2562), .CK(net_16632), .RN(x6501) );
DFFR_X2 inst_7193 ( .QN(net_8960), .D(net_2455), .CK(net_16153), .RN(x6501) );
CLKBUF_X2 inst_15347 ( .A(net_15194), .Z(net_15195) );
NAND2_X2 inst_4877 ( .A1(net_6152), .ZN(net_803), .A2(net_533) );
INV_X4 inst_5420 ( .ZN(net_1484), .A(net_858) );
CLKBUF_X2 inst_9994 ( .A(net_9841), .Z(net_9842) );
XOR2_X1 inst_94 ( .Z(net_1406), .B(net_1405), .A(net_610) );
CLKBUF_X2 inst_10946 ( .A(net_10793), .Z(net_10794) );
CLKBUF_X2 inst_18489 ( .A(net_18336), .Z(net_18337) );
CLKBUF_X2 inst_14615 ( .A(net_14462), .Z(net_14463) );
CLKBUF_X2 inst_17314 ( .A(net_17161), .Z(net_17162) );
CLKBUF_X2 inst_11858 ( .A(net_11705), .Z(net_11706) );
CLKBUF_X2 inst_13060 ( .A(net_12907), .Z(net_12908) );
SDFF_X2 inst_591 ( .SI(net_8382), .Q(net_8382), .SE(net_3969), .D(net_3962), .CK(net_12979) );
SDFF_X2 inst_424 ( .Q(net_8741), .D(net_8741), .SE(net_3982), .SI(net_3961), .CK(net_10199) );
NAND2_X2 inst_4345 ( .A1(net_7106), .A2(net_5164), .ZN(net_5112) );
CLKBUF_X2 inst_15504 ( .A(net_15351), .Z(net_15352) );
CLKBUF_X2 inst_15338 ( .A(net_14631), .Z(net_15186) );
CLKBUF_X2 inst_18721 ( .A(net_14232), .Z(net_18569) );
CLKBUF_X2 inst_10428 ( .A(net_10275), .Z(net_10276) );
CLKBUF_X2 inst_17624 ( .A(net_17471), .Z(net_17472) );
NAND2_X2 inst_4417 ( .A1(net_6856), .A2(net_5016), .ZN(net_5010) );
CLKBUF_X2 inst_10784 ( .A(net_10083), .Z(net_10632) );
AOI22_X2 inst_8320 ( .B1(net_8586), .A1(net_8475), .A2(net_6263), .B2(net_6262), .ZN(net_3726) );
INV_X4 inst_5727 ( .A(net_7626), .ZN(net_565) );
CLKBUF_X2 inst_14012 ( .A(net_9511), .Z(net_13860) );
CLKBUF_X2 inst_11861 ( .A(net_10114), .Z(net_11709) );
DFF_X1 inst_6853 ( .Q(net_6441), .D(net_3629), .CK(net_17956) );
SDFFR_X1 inst_2706 ( .QN(net_6799), .SE(net_6268), .SI(net_4360), .D(net_1235), .CK(net_11797), .RN(x6501) );
SDFF_X2 inst_476 ( .SI(net_8449), .Q(net_8449), .SE(net_3983), .D(net_3938), .CK(net_12469) );
AOI222_X1 inst_8640 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3933), .B1(net_3171), .C1(net_3170), .A1(x13772) );
CLKBUF_X2 inst_16389 ( .A(net_16236), .Z(net_16237) );
NAND4_X2 inst_3742 ( .ZN(net_4288), .A1(net_4064), .A2(net_4063), .A3(net_4062), .A4(net_4061) );
HA_X1 inst_6684 ( .A(net_3203), .S(net_3013), .CO(net_3012), .B(net_2971) );
CLKBUF_X2 inst_10249 ( .A(net_10096), .Z(net_10097) );
SDFFR_X2 inst_2499 ( .Q(net_8978), .D(net_8978), .SI(net_2618), .SE(net_2562), .CK(net_16636), .RN(x6501) );
CLKBUF_X2 inst_16150 ( .A(net_15997), .Z(net_15998) );
XOR2_X2 inst_20 ( .Z(net_1410), .B(net_1409), .A(net_615) );
CLKBUF_X2 inst_11542 ( .A(net_11389), .Z(net_11390) );
CLKBUF_X2 inst_18222 ( .A(net_18069), .Z(net_18070) );
CLKBUF_X2 inst_10007 ( .A(net_9134), .Z(net_9855) );
INV_X4 inst_5549 ( .ZN(net_813), .A(net_759) );
CLKBUF_X2 inst_13421 ( .A(net_9173), .Z(net_13269) );
MUX2_X2 inst_4994 ( .A(net_9021), .Z(net_3947), .B(net_1763), .S(net_622) );
CLKBUF_X2 inst_15387 ( .A(net_15234), .Z(net_15235) );
SDFF_X2 inst_576 ( .Q(net_8842), .D(net_8842), .SE(net_3964), .SI(net_3941), .CK(net_13423) );
CLKBUF_X2 inst_13590 ( .A(net_13437), .Z(net_13438) );
CLKBUF_X2 inst_14477 ( .A(net_14324), .Z(net_14325) );
CLKBUF_X2 inst_14398 ( .A(net_10602), .Z(net_14246) );
CLKBUF_X2 inst_10131 ( .A(net_9930), .Z(net_9979) );
CLKBUF_X2 inst_10182 ( .A(net_10029), .Z(net_10030) );
CLKBUF_X2 inst_17970 ( .A(net_17817), .Z(net_17818) );
CLKBUF_X2 inst_10376 ( .A(net_10223), .Z(net_10224) );
CLKBUF_X2 inst_16629 ( .A(net_16476), .Z(net_16477) );
OAI21_X2 inst_3055 ( .B2(net_8237), .B1(net_4850), .ZN(net_4755), .A(net_2607) );
OR2_X2 inst_2876 ( .ZN(net_4411), .A2(net_4406), .A1(net_4389) );
CLKBUF_X2 inst_16371 ( .A(net_16218), .Z(net_16219) );
CLKBUF_X2 inst_16516 ( .A(net_16363), .Z(net_16364) );
SDFF_X2 inst_976 ( .SI(net_7340), .Q(net_6747), .D(net_6747), .SE(net_3124), .CK(net_11911) );
CLKBUF_X2 inst_17150 ( .A(net_16997), .Z(net_16998) );
CLKBUF_X2 inst_9919 ( .A(net_9766), .Z(net_9767) );
CLKBUF_X2 inst_17610 ( .A(net_17457), .Z(net_17458) );
SDFF_X2 inst_1279 ( .Q(net_7838), .D(net_7838), .SE(net_2730), .SI(net_2656), .CK(net_16726) );
DFFR_X2 inst_7027 ( .QN(net_6292), .D(net_5683), .CK(net_16733), .RN(x6501) );
INV_X2 inst_6562 ( .A(net_9011), .ZN(net_492) );
CLKBUF_X2 inst_16437 ( .A(net_16284), .Z(net_16285) );
CLKBUF_X2 inst_16554 ( .A(net_11197), .Z(net_16402) );
DFFR_X1 inst_7474 ( .QN(net_7437), .D(net_4214), .CK(net_10118), .RN(x6501) );
CLKBUF_X2 inst_13011 ( .A(net_12858), .Z(net_12859) );
CLKBUF_X2 inst_13280 ( .A(net_13127), .Z(net_13128) );
CLKBUF_X2 inst_13287 ( .A(net_13134), .Z(net_13135) );
AOI22_X2 inst_8025 ( .B1(net_8134), .A1(net_7896), .A2(net_6098), .B2(net_4190), .ZN(net_4112) );
CLKBUF_X2 inst_11036 ( .A(net_10883), .Z(net_10884) );
CLKBUF_X2 inst_18145 ( .A(net_17992), .Z(net_17993) );
NOR2_X2 inst_3414 ( .A1(net_8898), .ZN(net_3362), .A2(net_3151) );
NOR2_X2 inst_3399 ( .ZN(net_4358), .A2(net_4357), .A1(net_704) );
CLKBUF_X2 inst_17223 ( .A(net_14343), .Z(net_17071) );
NAND2_X2 inst_4495 ( .ZN(net_4477), .A2(net_4388), .A1(net_2602) );
SDFF_X2 inst_1432 ( .SI(net_7272), .Q(net_7049), .D(net_7049), .SE(net_6280), .CK(net_16856) );
INV_X4 inst_5667 ( .A(net_6351), .ZN(net_579) );
CLKBUF_X2 inst_12159 ( .A(net_10313), .Z(net_12007) );
OAI21_X2 inst_3084 ( .ZN(net_3179), .A(net_2998), .B2(net_2996), .B1(net_1206) );
CLKBUF_X2 inst_19006 ( .A(net_18853), .Z(net_18854) );
CLKBUF_X2 inst_11739 ( .A(net_11586), .Z(net_11587) );
CLKBUF_X2 inst_15562 ( .A(net_15409), .Z(net_15410) );
CLKBUF_X2 inst_16344 ( .A(net_16191), .Z(net_16192) );
SDFFR_X2 inst_2464 ( .SE(net_2260), .Q(net_328), .D(net_328), .CK(net_10399), .RN(x6501), .SI(x2746) );
CLKBUF_X2 inst_9790 ( .A(net_9637), .Z(net_9638) );
AOI221_X2 inst_8776 ( .B2(net_8238), .B1(net_5268), .C2(net_5267), .ZN(net_5263), .A(net_4913), .C1(net_175) );
CLKBUF_X2 inst_9433 ( .A(net_9280), .Z(net_9281) );
CLKBUF_X2 inst_11197 ( .A(net_11044), .Z(net_11045) );
CLKBUF_X2 inst_14432 ( .A(net_11348), .Z(net_14280) );
CLKBUF_X2 inst_16347 ( .A(net_16194), .Z(net_16195) );
NAND3_X2 inst_4010 ( .ZN(net_1910), .A2(net_1085), .A1(net_1060), .A3(net_686) );
CLKBUF_X2 inst_15373 ( .A(net_15220), .Z(net_15221) );
NOR2_X4 inst_3328 ( .ZN(net_3359), .A1(net_3160), .A2(net_3074) );
CLKBUF_X2 inst_9677 ( .A(net_9524), .Z(net_9525) );
CLKBUF_X2 inst_13254 ( .A(net_13101), .Z(net_13102) );
AOI22_X2 inst_8399 ( .B1(net_8711), .A1(net_8489), .B2(net_4350), .A2(net_4349), .ZN(net_3653) );
SDFF_X2 inst_1111 ( .D(net_7342), .SI(net_6551), .Q(net_6551), .SE(net_3086), .CK(net_9459) );
CLKBUF_X2 inst_14495 ( .A(net_14342), .Z(net_14343) );
CLKBUF_X2 inst_17925 ( .A(net_16284), .Z(net_17773) );
SDFFR_X1 inst_2658 ( .D(net_6780), .SE(net_4506), .CK(net_11416), .RN(x6501), .SI(x1467), .Q(x1467) );
AND2_X4 inst_9122 ( .A2(net_6753), .A1(net_6752), .ZN(net_2902) );
CLKBUF_X2 inst_11496 ( .A(net_11343), .Z(net_11344) );
SDFF_X2 inst_480 ( .SI(net_8454), .Q(net_8454), .SE(net_3983), .D(net_3946), .CK(net_11100) );
NAND2_X2 inst_4631 ( .ZN(net_2514), .A1(net_2473), .A2(net_2404) );
OAI21_X2 inst_2986 ( .ZN(net_5913), .B2(net_5912), .A(net_5804), .B1(net_702) );
SDFFR_X2 inst_2206 ( .SI(net_8941), .Q(net_8941), .SE(net_6144), .D(net_1609), .CK(net_16261), .RN(x6501) );
AOI22_X2 inst_8074 ( .B1(net_8073), .A1(net_7869), .B2(net_6107), .A2(net_4400), .ZN(net_4070) );
OR4_X4 inst_2792 ( .A1(net_7616), .A4(net_6180), .A3(net_5691), .ZN(net_3093), .A2(net_2429) );
CLKBUF_X2 inst_13597 ( .A(net_13341), .Z(net_13445) );
CLKBUF_X2 inst_17053 ( .A(net_16900), .Z(net_16901) );
SDFF_X2 inst_739 ( .Q(net_8812), .D(net_8812), .SI(net_3939), .SE(net_3879), .CK(net_12526) );
CLKBUF_X2 inst_18111 ( .A(net_17400), .Z(net_17959) );
XOR2_X2 inst_46 ( .A(net_1763), .Z(net_1019), .B(net_593) );
INV_X16 inst_6637 ( .ZN(net_3979), .A(net_3353) );
SDFFR_X2 inst_2537 ( .QN(net_6374), .SE(net_2147), .SI(net_1951), .D(net_683), .CK(net_14956), .RN(x6501) );
CLKBUF_X2 inst_15530 ( .A(net_15377), .Z(net_15378) );
CLKBUF_X2 inst_16862 ( .A(net_16709), .Z(net_16710) );
SDFF_X2 inst_1126 ( .D(net_7332), .SI(net_6574), .Q(net_6574), .SE(net_3070), .CK(net_9416) );
CLKBUF_X2 inst_12361 ( .A(net_9701), .Z(net_12209) );
CLKBUF_X2 inst_16180 ( .A(net_14614), .Z(net_16028) );
NOR2_X2 inst_3470 ( .ZN(net_2449), .A1(net_2349), .A2(net_2297) );
CLKBUF_X2 inst_13065 ( .A(net_9304), .Z(net_12913) );
SDFF_X2 inst_796 ( .SI(net_8368), .Q(net_8368), .D(net_3939), .SE(net_3880), .CK(net_10514) );
CLKBUF_X2 inst_14135 ( .A(net_13982), .Z(net_13983) );
CLKBUF_X2 inst_16253 ( .A(net_16100), .Z(net_16101) );
CLKBUF_X2 inst_11727 ( .A(net_11574), .Z(net_11575) );
HA_X1 inst_6699 ( .S(net_2564), .CO(net_2563), .B(net_2390), .A(x3288) );
CLKBUF_X2 inst_15030 ( .A(net_12913), .Z(net_14878) );
SDFF_X2 inst_1499 ( .SI(net_7857), .Q(net_7857), .D(net_2719), .SE(net_2558), .CK(net_18795) );
OAI221_X2 inst_2972 ( .B2(net_2489), .C2(net_2450), .ZN(net_2422), .A(net_2272), .B1(net_1272), .C1(net_659) );
CLKBUF_X2 inst_9470 ( .A(net_9071), .Z(net_9318) );
CLKBUF_X2 inst_15554 ( .A(net_15401), .Z(net_15402) );
CLKBUF_X2 inst_9293 ( .A(net_9140), .Z(net_9141) );
CLKBUF_X2 inst_12345 ( .A(net_12192), .Z(net_12193) );
NOR3_X2 inst_3297 ( .A1(net_6159), .ZN(net_4728), .A2(net_1887), .A3(net_1886) );
INV_X4 inst_5931 ( .A(net_7307), .ZN(net_1236) );
INV_X4 inst_5429 ( .A(net_1267), .ZN(net_1104) );
CLKBUF_X2 inst_18823 ( .A(net_18670), .Z(net_18671) );
CLKBUF_X2 inst_12556 ( .A(net_12403), .Z(net_12404) );
NAND2_X2 inst_4423 ( .A1(net_6861), .A2(net_5016), .ZN(net_5004) );
CLKBUF_X2 inst_10438 ( .A(net_10285), .Z(net_10286) );
CLKBUF_X2 inst_13384 ( .A(net_13231), .Z(net_13232) );
CLKBUF_X2 inst_11880 ( .A(net_11727), .Z(net_11728) );
NAND2_X2 inst_4342 ( .A1(net_7105), .A2(net_5164), .ZN(net_5115) );
CLKBUF_X2 inst_15691 ( .A(net_15538), .Z(net_15539) );
AOI222_X1 inst_8664 ( .A2(net_3599), .B2(net_3598), .C2(net_3597), .ZN(net_3594), .C1(net_3082), .A1(net_1568), .B1(net_1452) );
CLKBUF_X2 inst_10398 ( .A(net_10245), .Z(net_10246) );
CLKBUF_X2 inst_12887 ( .A(net_12734), .Z(net_12735) );
NAND2_X2 inst_4339 ( .A1(net_7104), .A2(net_5164), .ZN(net_5118) );
INV_X8 inst_5060 ( .ZN(net_6273), .A(net_6272) );
CLKBUF_X2 inst_17666 ( .A(net_9344), .Z(net_17514) );
CLKBUF_X2 inst_14187 ( .A(net_11375), .Z(net_14035) );
SDFF_X2 inst_1421 ( .SI(net_7274), .Q(net_7051), .D(net_7051), .SE(net_6280), .CK(net_14144) );
CLKBUF_X2 inst_18909 ( .A(net_18756), .Z(net_18757) );
CLKBUF_X2 inst_16836 ( .A(net_16643), .Z(net_16684) );
NAND2_X2 inst_4262 ( .A1(net_7033), .A2(net_5249), .ZN(net_5198) );
CLKBUF_X2 inst_12819 ( .A(net_12666), .Z(net_12667) );
AOI22_X2 inst_8298 ( .B1(net_8806), .A1(net_8547), .ZN(net_6230), .A2(net_3861), .B2(net_3860) );
CLKBUF_X2 inst_12607 ( .A(net_11540), .Z(net_12455) );
CLKBUF_X2 inst_10406 ( .A(net_9576), .Z(net_10254) );
CLKBUF_X2 inst_16283 ( .A(net_16130), .Z(net_16131) );
CLKBUF_X2 inst_17797 ( .A(net_17644), .Z(net_17645) );
CLKBUF_X2 inst_17436 ( .A(net_17283), .Z(net_17284) );
CLKBUF_X2 inst_13882 ( .A(net_13729), .Z(net_13730) );
NAND4_X2 inst_3664 ( .A4(net_6018), .A1(net_6017), .ZN(net_4601), .A2(net_4108), .A3(net_4107) );
CLKBUF_X2 inst_9688 ( .A(net_9535), .Z(net_9536) );
CLKBUF_X2 inst_9961 ( .A(net_9415), .Z(net_9809) );
INV_X4 inst_6011 ( .A(net_6369), .ZN(net_933) );
CLKBUF_X2 inst_10536 ( .A(net_9063), .Z(net_10384) );
CLKBUF_X2 inst_18437 ( .A(net_18284), .Z(net_18285) );
CLKBUF_X2 inst_17412 ( .A(net_17259), .Z(net_17260) );
NOR2_X2 inst_3486 ( .A1(net_2290), .ZN(net_2119), .A2(net_1917) );
AOI221_X2 inst_8833 ( .C1(net_8168), .B1(net_7726), .C2(net_6101), .B2(net_6095), .ZN(net_6015), .A(net_4296) );
CLKBUF_X2 inst_13246 ( .A(net_13093), .Z(net_13094) );
CLKBUF_X2 inst_13961 ( .A(net_13808), .Z(net_13809) );
CLKBUF_X2 inst_9636 ( .A(net_9483), .Z(net_9484) );
AOI21_X2 inst_8970 ( .B2(net_5947), .ZN(net_2588), .A(net_2587), .B1(net_916) );
CLKBUF_X2 inst_12099 ( .A(net_10934), .Z(net_11947) );
CLKBUF_X2 inst_13358 ( .A(net_11194), .Z(net_13206) );
CLKBUF_X2 inst_13769 ( .A(net_9063), .Z(net_13617) );
CLKBUF_X2 inst_18987 ( .A(net_14432), .Z(net_18835) );
INV_X16 inst_6628 ( .ZN(net_3860), .A(net_3383) );
CLKBUF_X2 inst_17257 ( .A(net_17104), .Z(net_17105) );
CLKBUF_X2 inst_10029 ( .A(net_9681), .Z(net_9877) );
CLKBUF_X2 inst_13877 ( .A(net_13724), .Z(net_13725) );
XNOR2_X2 inst_230 ( .B(net_4890), .ZN(net_1312), .A(net_1099) );
INV_X4 inst_5903 ( .A(net_6303), .ZN(net_2687) );
CLKBUF_X2 inst_18022 ( .A(net_17869), .Z(net_17870) );
CLKBUF_X2 inst_18982 ( .A(net_18829), .Z(net_18830) );
CLKBUF_X2 inst_16668 ( .A(net_16515), .Z(net_16516) );
CLKBUF_X2 inst_10089 ( .A(net_9936), .Z(net_9937) );
CLKBUF_X2 inst_17337 ( .A(net_17184), .Z(net_17185) );
SDFF_X2 inst_1893 ( .D(net_7278), .SI(net_7015), .Q(net_7015), .SE(net_6277), .CK(net_14610) );
INV_X4 inst_5101 ( .ZN(net_5692), .A(net_5660) );
NAND2_X2 inst_4728 ( .ZN(net_2658), .A2(net_1586), .A1(net_1225) );
CLKBUF_X2 inst_16074 ( .A(net_13761), .Z(net_15922) );
INV_X2 inst_6480 ( .ZN(net_907), .A(net_230) );
AOI22_X2 inst_8325 ( .A1(net_8623), .B1(net_8438), .A2(net_3864), .B2(net_3863), .ZN(net_3721) );
NAND2_X2 inst_4385 ( .A1(net_7078), .A2(net_5162), .ZN(net_5072) );
CLKBUF_X2 inst_16841 ( .A(net_12508), .Z(net_16689) );
NAND2_X2 inst_4606 ( .A2(net_6144), .ZN(net_2629), .A1(net_2628) );
CLKBUF_X2 inst_18986 ( .A(net_10910), .Z(net_18834) );
CLKBUF_X2 inst_17782 ( .A(net_17629), .Z(net_17630) );
CLKBUF_X2 inst_18472 ( .A(net_18319), .Z(net_18320) );
SDFF_X2 inst_452 ( .Q(net_8750), .D(net_8750), .SE(net_3982), .SI(net_3946), .CK(net_10769) );
CLKBUF_X2 inst_14375 ( .A(net_14222), .Z(net_14223) );
CLKBUF_X2 inst_18603 ( .A(net_18450), .Z(net_18451) );
CLKBUF_X2 inst_17088 ( .A(net_16935), .Z(net_16936) );
CLKBUF_X2 inst_10338 ( .A(net_10185), .Z(net_10186) );
CLKBUF_X2 inst_9392 ( .A(net_9239), .Z(net_9240) );
AOI22_X2 inst_8397 ( .B1(net_8563), .A1(net_8452), .A2(net_6263), .B2(net_6262), .ZN(net_3655) );
OAI21_X2 inst_3061 ( .B2(net_8245), .B1(net_4850), .ZN(net_4746), .A(net_2601) );
CLKBUF_X2 inst_13146 ( .A(net_12993), .Z(net_12994) );
NAND2_X2 inst_4144 ( .ZN(net_5375), .A2(net_5214), .A1(net_5111) );
CLKBUF_X2 inst_14000 ( .A(net_13847), .Z(net_13848) );
CLKBUF_X2 inst_17953 ( .A(net_14769), .Z(net_17801) );
CLKBUF_X2 inst_17710 ( .A(net_17557), .Z(net_17558) );
CLKBUF_X2 inst_10254 ( .A(net_9196), .Z(net_10102) );
SDFF_X2 inst_728 ( .SI(net_8494), .Q(net_8494), .D(net_3945), .SE(net_3884), .CK(net_13099) );
CLKBUF_X2 inst_11180 ( .A(net_11027), .Z(net_11028) );
CLKBUF_X2 inst_14308 ( .A(net_9842), .Z(net_14156) );
CLKBUF_X2 inst_10372 ( .A(net_10219), .Z(net_10220) );
OAI21_X2 inst_3121 ( .ZN(net_2349), .A(net_2296), .B2(net_2290), .B1(net_149) );
SDFFR_X1 inst_2780 ( .Q(net_7283), .D(net_2803), .SI(net_1867), .SE(net_1327), .CK(net_18163), .RN(x6501) );
CLKBUF_X2 inst_15034 ( .A(net_14881), .Z(net_14882) );
INV_X1 inst_6655 ( .A(net_6155), .ZN(net_6153) );
CLKBUF_X2 inst_18957 ( .A(net_18804), .Z(net_18805) );
NAND2_X2 inst_4152 ( .ZN(net_5364), .A1(net_5104), .A2(net_5103) );
CLKBUF_X2 inst_16325 ( .A(net_12241), .Z(net_16173) );
CLKBUF_X2 inst_11031 ( .A(net_10878), .Z(net_10879) );
OR2_X4 inst_2844 ( .A2(net_3262), .ZN(net_1880), .A1(net_1787) );
CLKBUF_X2 inst_19178 ( .A(net_17429), .Z(net_19026) );
SDFFR_X2 inst_2492 ( .Q(net_8987), .D(net_8987), .SI(net_2592), .SE(net_2562), .CK(net_16407), .RN(x6501) );
CLKBUF_X2 inst_17046 ( .A(net_16893), .Z(net_16894) );
NOR2_X2 inst_3582 ( .A2(net_7524), .A1(net_1480), .ZN(net_1372) );
CLKBUF_X2 inst_15571 ( .A(net_13371), .Z(net_15419) );
NOR2_X2 inst_3480 ( .ZN(net_2402), .A1(net_2244), .A2(net_2076) );
CLKBUF_X2 inst_14125 ( .A(net_13972), .Z(net_13973) );
CLKBUF_X2 inst_18114 ( .A(net_17961), .Z(net_17962) );
CLKBUF_X2 inst_11721 ( .A(net_11568), .Z(net_11569) );
INV_X4 inst_5705 ( .ZN(net_2555), .A(net_433) );
CLKBUF_X2 inst_10879 ( .A(net_10726), .Z(net_10727) );
CLKBUF_X2 inst_15314 ( .A(net_15161), .Z(net_15162) );
CLKBUF_X2 inst_14776 ( .A(net_12180), .Z(net_14624) );
DFFR_X2 inst_7093 ( .QN(net_7213), .D(net_3387), .CK(net_18963), .RN(x6501) );
CLKBUF_X2 inst_11017 ( .A(net_10864), .Z(net_10865) );
NAND2_X2 inst_4818 ( .ZN(net_1246), .A1(net_896), .A2(net_611) );
CLKBUF_X2 inst_10381 ( .A(net_10228), .Z(net_10229) );
SDFF_X2 inst_974 ( .SI(net_7337), .Q(net_6744), .D(net_6744), .SE(net_3124), .CK(net_9504) );
CLKBUF_X2 inst_17685 ( .A(net_17532), .Z(net_17533) );
CLKBUF_X2 inst_18700 ( .A(net_18547), .Z(net_18548) );
SDFF_X2 inst_1001 ( .D(net_7341), .SI(net_6649), .Q(net_6649), .SE(net_3123), .CK(net_9494) );
CLKBUF_X2 inst_17281 ( .A(net_17128), .Z(net_17129) );
INV_X4 inst_5825 ( .ZN(net_2800), .A(net_266) );
OAI21_X2 inst_3033 ( .ZN(net_4851), .B1(net_4850), .B2(net_4849), .A(net_2619) );
OAI22_X2 inst_2925 ( .A2(net_2967), .B2(net_2943), .ZN(net_2893), .A1(net_1533), .B1(net_1135) );
AOI22_X2 inst_7843 ( .A2(net_5595), .ZN(net_4665), .B2(net_4388), .B1(net_2618), .A1(net_313) );
CLKBUF_X2 inst_10537 ( .A(net_10384), .Z(net_10385) );
SDFF_X2 inst_1828 ( .D(net_7285), .SI(net_6862), .Q(net_6862), .SE(net_6282), .CK(net_16195) );
CLKBUF_X2 inst_9510 ( .A(net_9357), .Z(net_9358) );
NOR2_X2 inst_3388 ( .A1(net_4898), .ZN(net_4779), .A2(net_4640) );
NAND4_X2 inst_3735 ( .ZN(net_4295), .A1(net_4106), .A2(net_4105), .A3(net_4104), .A4(net_4103) );
CLKBUF_X2 inst_11238 ( .A(net_9685), .Z(net_11086) );
INV_X4 inst_5311 ( .A(net_1607), .ZN(net_1474) );
SDFFR_X1 inst_2675 ( .SI(net_7537), .SE(net_5043), .CK(net_9712), .RN(x6501), .Q(x4093), .D(x4093) );
CLKBUF_X2 inst_18115 ( .A(net_12230), .Z(net_17963) );
XNOR2_X2 inst_141 ( .A(net_2433), .ZN(net_2326), .B(net_2277) );
SDFFR_X2 inst_2520 ( .SI(net_7217), .Q(net_7217), .D(net_2167), .SE(net_1379), .CK(net_18907), .RN(x6501) );
CLKBUF_X2 inst_10578 ( .A(net_10425), .Z(net_10426) );
SDFF_X2 inst_571 ( .Q(net_8835), .D(net_8835), .SE(net_3964), .SI(net_3957), .CK(net_12337) );
CLKBUF_X2 inst_16405 ( .A(net_16252), .Z(net_16253) );
INV_X4 inst_6007 ( .A(net_7592), .ZN(net_511) );
SDFF_X2 inst_1974 ( .D(net_7302), .SI(net_6919), .Q(net_6919), .SE(net_6284), .CK(net_15395) );
SDFF_X2 inst_2017 ( .SI(net_7799), .Q(net_7799), .D(net_2639), .SE(net_2459), .CK(net_14381) );
SDFF_X2 inst_1154 ( .SI(net_7336), .Q(net_6611), .D(net_6611), .SE(net_3069), .CK(net_9449) );
CLKBUF_X2 inst_14901 ( .A(net_11128), .Z(net_14749) );
CLKBUF_X2 inst_16267 ( .A(net_16114), .Z(net_16115) );
CLKBUF_X1 inst_7728 ( .A(x192486), .Z(x1010) );
CLKBUF_X2 inst_12413 ( .A(net_11574), .Z(net_12261) );
CLKBUF_X2 inst_9584 ( .A(net_9431), .Z(net_9432) );
CLKBUF_X2 inst_16339 ( .A(net_16186), .Z(net_16187) );
DFFR_X2 inst_7224 ( .QN(net_8962), .D(net_2237), .CK(net_14480), .RN(x6501) );
SDFF_X2 inst_469 ( .SI(net_8447), .Q(net_8447), .SE(net_3983), .D(net_3980), .CK(net_13359) );
DFFR_X1 inst_7468 ( .QN(net_7432), .D(net_4271), .CK(net_12398), .RN(x6501) );
AOI222_X1 inst_8598 ( .B2(net_6777), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5827), .A1(net_3043), .C1(x2693) );
DFFR_X2 inst_7133 ( .QN(net_7637), .D(net_3034), .CK(net_18953), .RN(x6501) );
DFF_X1 inst_6837 ( .QN(net_6456), .D(net_3611), .CK(net_17908) );
CLKBUF_X2 inst_15013 ( .A(net_14860), .Z(net_14861) );
CLKBUF_X2 inst_16919 ( .A(net_16766), .Z(net_16767) );
AOI21_X4 inst_8866 ( .A(net_6254), .ZN(net_5934), .B2(net_5918), .B1(net_4372) );
INV_X16 inst_6642 ( .ZN(net_4345), .A(net_3316) );
INV_X2 inst_6507 ( .A(net_7578), .ZN(net_3140) );
SDFFR_X2 inst_2339 ( .D(net_7372), .SI(net_2737), .SE(net_2734), .QN(net_275), .CK(net_14555), .RN(x6501) );
CLKBUF_X2 inst_18911 ( .A(net_16125), .Z(net_18759) );
CLKBUF_X2 inst_12300 ( .A(net_12147), .Z(net_12148) );
CLKBUF_X2 inst_18692 ( .A(net_18539), .Z(net_18540) );
CLKBUF_X2 inst_11603 ( .A(net_9914), .Z(net_11451) );
SDFF_X2 inst_1216 ( .Q(net_7963), .D(net_7963), .SE(net_2755), .SI(net_2713), .CK(net_14299) );
AOI22_X2 inst_8260 ( .B1(net_8578), .A1(net_8467), .A2(net_6263), .B2(net_6262), .ZN(net_3778) );
HA_X1 inst_6697 ( .B(net_6136), .A(net_2916), .S(net_2568), .CO(net_2567) );
CLKBUF_X2 inst_15544 ( .A(net_15391), .Z(net_15392) );
CLKBUF_X2 inst_17019 ( .A(net_11976), .Z(net_16867) );
SDFF_X2 inst_952 ( .SI(net_7338), .Q(net_6712), .D(net_6712), .SE(net_3125), .CK(net_9506) );
CLKBUF_X2 inst_18833 ( .A(net_18680), .Z(net_18681) );
CLKBUF_X2 inst_16069 ( .A(net_13628), .Z(net_15917) );
INV_X4 inst_5972 ( .A(net_7621), .ZN(net_1563) );
DFFR_X2 inst_7254 ( .QN(net_7398), .D(net_1969), .CK(net_17866), .RN(x6501) );
CLKBUF_X2 inst_14710 ( .A(net_14557), .Z(net_14558) );
SDFF_X2 inst_721 ( .SI(net_8505), .Q(net_8505), .D(net_3942), .SE(net_3884), .CK(net_12593) );
CLKBUF_X2 inst_11135 ( .A(net_10982), .Z(net_10983) );
DFFR_X2 inst_7211 ( .D(net_2362), .QN(net_216), .CK(net_17469), .RN(x6501) );
CLKBUF_X2 inst_10838 ( .A(net_10685), .Z(net_10686) );
OAI21_X2 inst_3009 ( .B2(net_5755), .ZN(net_5723), .A(net_5719), .B1(net_494) );
SDFF_X2 inst_1366 ( .Q(net_8015), .D(net_8015), .SI(net_2659), .SE(net_2545), .CK(net_15533) );
CLKBUF_X2 inst_13667 ( .A(net_13514), .Z(net_13515) );
CLKBUF_X2 inst_13079 ( .A(net_9666), .Z(net_12927) );
CLKBUF_X2 inst_17675 ( .A(net_17522), .Z(net_17523) );
SDFF_X2 inst_1915 ( .D(net_7289), .SI(net_6906), .Q(net_6906), .SE(net_6284), .CK(net_15311) );
OR4_X2 inst_2794 ( .A3(net_8941), .A1(net_2680), .ZN(net_2409), .A2(net_2408), .A4(net_2221) );
SDFF_X2 inst_1254 ( .SI(net_7676), .Q(net_7676), .SE(net_2714), .D(net_2708), .CK(net_18294) );
DFFR_X2 inst_7111 ( .QN(net_8258), .D(net_3220), .CK(net_18500), .RN(x6501) );
NOR2_X2 inst_3553 ( .ZN(net_4324), .A2(net_4320), .A1(net_1380) );
CLKBUF_X2 inst_14031 ( .A(net_11624), .Z(net_13879) );
CLKBUF_X2 inst_14412 ( .A(net_14259), .Z(net_14260) );
SDFF_X2 inst_1811 ( .SI(net_8057), .Q(net_8057), .D(net_2720), .SE(net_2508), .CK(net_18032) );
NAND2_X2 inst_4544 ( .A2(net_3356), .ZN(net_3350), .A1(net_3318) );
CLKBUF_X2 inst_11147 ( .A(net_10994), .Z(net_10995) );
CLKBUF_X2 inst_11351 ( .A(net_10523), .Z(net_11199) );
CLKBUF_X2 inst_14479 ( .A(net_14326), .Z(net_14327) );
CLKBUF_X2 inst_10801 ( .A(net_10648), .Z(net_10649) );
DFFR_X2 inst_7054 ( .QN(net_7507), .D(net_4786), .CK(net_14833), .RN(x6501) );
CLKBUF_X2 inst_18075 ( .A(net_11184), .Z(net_17923) );
CLKBUF_X2 inst_14834 ( .A(net_14681), .Z(net_14682) );
AOI221_X2 inst_8826 ( .B1(net_8056), .C1(net_7852), .B2(net_6107), .ZN(net_5999), .C2(net_4400), .A(net_4307) );
XNOR2_X2 inst_163 ( .ZN(net_1844), .A(net_1487), .B(net_662) );
AND2_X2 inst_9156 ( .ZN(net_2865), .A2(net_2864), .A1(net_2661) );
SDFF_X2 inst_394 ( .Q(net_8830), .D(net_8830), .SI(net_3973), .SE(net_3964), .CK(net_13216) );
AOI22_X2 inst_8455 ( .B1(net_6604), .A1(net_6571), .A2(net_6257), .B2(net_6110), .ZN(net_3485) );
CLKBUF_X2 inst_11619 ( .A(net_9413), .Z(net_11467) );
CLKBUF_X2 inst_18978 ( .A(net_18101), .Z(net_18826) );
CLKBUF_X2 inst_17678 ( .A(net_17525), .Z(net_17526) );
CLKBUF_X2 inst_16268 ( .A(net_9537), .Z(net_16116) );
SDFF_X2 inst_1814 ( .D(net_7281), .SI(net_7018), .Q(net_7018), .SE(net_6277), .CK(net_19007) );
NAND2_X2 inst_4470 ( .A1(net_5588), .ZN(net_4704), .A2(net_4642) );
CLKBUF_X2 inst_17392 ( .A(net_17239), .Z(net_17240) );
CLKBUF_X2 inst_10875 ( .A(net_9545), .Z(net_10723) );
SDFF_X2 inst_361 ( .Q(net_8752), .D(net_8752), .SE(net_3982), .SI(net_3962), .CK(net_10208) );
CLKBUF_X2 inst_11358 ( .A(net_11205), .Z(net_11206) );
NOR2_X2 inst_3400 ( .A1(net_6197), .ZN(net_4403), .A2(net_4357) );
AOI22_X2 inst_8127 ( .B1(net_8083), .A1(net_7743), .B2(net_6108), .A2(net_6096), .ZN(net_4022) );
CLKBUF_X2 inst_12134 ( .A(net_11803), .Z(net_11982) );
AOI22_X2 inst_8082 ( .B1(net_8080), .A1(net_7740), .B2(net_6108), .A2(net_6096), .ZN(net_4063) );
CLKBUF_X2 inst_19056 ( .A(net_18903), .Z(net_18904) );
CLKBUF_X2 inst_11008 ( .A(net_10855), .Z(net_10856) );
CLKBUF_X2 inst_14852 ( .A(net_14699), .Z(net_14700) );
SDFF_X2 inst_786 ( .SI(net_8356), .Q(net_8356), .D(net_3963), .SE(net_3880), .CK(net_10901) );
XOR2_X2 inst_2 ( .Z(net_3218), .A(net_3042), .B(x2633) );
CLKBUF_X2 inst_11003 ( .A(net_10850), .Z(net_10851) );
SDFF_X2 inst_888 ( .Q(net_8559), .D(net_8559), .SI(net_3977), .SE(net_3878), .CK(net_11041) );
SDFF_X2 inst_1769 ( .D(net_7294), .SI(net_6871), .Q(net_6871), .SE(net_6282), .CK(net_17688) );
CLKBUF_X2 inst_12306 ( .A(net_12153), .Z(net_12154) );
INV_X4 inst_5999 ( .ZN(net_2697), .A(net_145) );
NAND4_X4 inst_3625 ( .ZN(net_2002), .A3(net_1646), .A2(net_1644), .A4(net_1554), .A1(net_1550) );
INV_X2 inst_6598 ( .A(net_6136), .ZN(net_6135) );
INV_X4 inst_5979 ( .ZN(net_2499), .A(net_231) );
CLKBUF_X2 inst_15896 ( .A(net_15743), .Z(net_15744) );
AOI22_X2 inst_7817 ( .A2(net_8226), .B2(net_6144), .A1(net_4764), .ZN(net_4737), .B1(net_4736) );
SDFFR_X2 inst_2581 ( .D(net_7385), .QN(net_7245), .SI(net_1955), .SE(net_1379), .CK(net_18114), .RN(x6501) );
NAND2_X2 inst_4110 ( .ZN(net_5420), .A1(net_5146), .A2(net_5145) );
SDFFR_X2 inst_2164 ( .QN(net_7585), .D(net_3955), .SE(net_3144), .SI(net_482), .CK(net_11032), .RN(x6501) );
CLKBUF_X2 inst_17112 ( .A(net_16959), .Z(net_16960) );
CLKBUF_X2 inst_16618 ( .A(net_16465), .Z(net_16466) );
DFFR_X2 inst_7198 ( .D(net_2361), .QN(net_217), .CK(net_17570), .RN(x6501) );
CLKBUF_X2 inst_13208 ( .A(net_13055), .Z(net_13056) );
NAND2_X2 inst_4392 ( .A1(net_7124), .A2(net_5166), .ZN(net_5065) );
CLKBUF_X2 inst_11696 ( .A(net_11543), .Z(net_11544) );
CLKBUF_X2 inst_11093 ( .A(net_10940), .Z(net_10941) );
MUX2_X2 inst_4915 ( .Z(net_5925), .S(net_5814), .B(net_5778), .A(net_3258) );
AOI222_X2 inst_8590 ( .B2(net_8246), .C1(net_7513), .A1(net_6214), .B1(net_4891), .C2(net_4889), .ZN(net_4804), .A2(net_4803) );
CLKBUF_X2 inst_14424 ( .A(net_14271), .Z(net_14272) );
CLKBUF_X2 inst_15758 ( .A(net_15605), .Z(net_15606) );
AOI22_X2 inst_8530 ( .B1(net_6657), .A1(net_6624), .A2(net_6213), .B2(net_6138), .ZN(net_3410) );
CLKBUF_X2 inst_9655 ( .A(net_9502), .Z(net_9503) );
CLKBUF_X2 inst_11245 ( .A(net_9689), .Z(net_11093) );
CLKBUF_X2 inst_16276 ( .A(net_16123), .Z(net_16124) );
CLKBUF_X2 inst_16926 ( .A(net_9643), .Z(net_16774) );
CLKBUF_X2 inst_17385 ( .A(net_14678), .Z(net_17233) );
NOR2_X2 inst_3385 ( .ZN(net_5466), .A2(net_5020), .A1(net_1787) );
SDFF_X2 inst_1572 ( .SI(net_7718), .Q(net_7718), .D(net_2589), .SE(net_2559), .CK(net_18386) );
CLKBUF_X2 inst_11753 ( .A(net_11600), .Z(net_11601) );
NAND2_X2 inst_4906 ( .A2(net_8950), .A1(net_8949), .ZN(net_1322) );
CLKBUF_X2 inst_16550 ( .A(net_9790), .Z(net_16398) );
CLKBUF_X2 inst_14932 ( .A(net_14779), .Z(net_14780) );
CLKBUF_X2 inst_14815 ( .A(net_14662), .Z(net_14663) );
CLKBUF_X2 inst_15634 ( .A(net_13393), .Z(net_15482) );
CLKBUF_X2 inst_14026 ( .A(net_13873), .Z(net_13874) );
CLKBUF_X2 inst_10221 ( .A(net_10068), .Z(net_10069) );
MUX2_X2 inst_4978 ( .A(net_9017), .Z(net_3980), .S(net_622), .B(net_569) );
CLKBUF_X2 inst_18608 ( .A(net_18455), .Z(net_18456) );
AOI22_X2 inst_7875 ( .A2(net_6440), .A1(net_5654), .B2(net_4881), .ZN(net_4566), .B1(net_240) );
CLKBUF_X2 inst_18787 ( .A(net_18634), .Z(net_18635) );
CLKBUF_X2 inst_9721 ( .A(net_9523), .Z(net_9569) );
CLKBUF_X2 inst_12048 ( .A(net_11895), .Z(net_11896) );
NAND2_X2 inst_4367 ( .A1(net_7072), .A2(net_5162), .ZN(net_5090) );
CLKBUF_X2 inst_10346 ( .A(net_10193), .Z(net_10194) );
SDFF_X2 inst_1731 ( .SI(net_7741), .Q(net_7741), .D(net_2655), .SE(net_2560), .CK(net_15481) );
CLKBUF_X2 inst_16631 ( .A(net_16478), .Z(net_16479) );
AOI22_X2 inst_7960 ( .B1(net_7922), .A1(net_7820), .B2(net_6103), .A2(net_4398), .ZN(net_4168) );
OAI221_X2 inst_2960 ( .ZN(net_4638), .B2(net_4553), .B1(net_4510), .C1(net_2981), .A(net_2939), .C2(net_1627) );
SDFF_X2 inst_1909 ( .D(net_7278), .SI(net_6975), .Q(net_6975), .SE(net_6283), .CK(net_14605) );
CLKBUF_X2 inst_16674 ( .A(net_16521), .Z(net_16522) );
INV_X2 inst_6616 ( .A(net_6211), .ZN(net_6210) );
NAND2_X2 inst_4318 ( .A1(net_7098), .A2(net_5164), .ZN(net_5139) );
CLKBUF_X2 inst_11080 ( .A(net_10927), .Z(net_10928) );
CLKBUF_X2 inst_11669 ( .A(net_11516), .Z(net_11517) );
AOI22_X2 inst_7991 ( .B1(net_7926), .A1(net_7824), .B2(net_6103), .A2(net_4398), .ZN(net_4141) );
AND2_X4 inst_9063 ( .ZN(net_6213), .A2(net_3250), .A1(net_3247) );
DFFR_X1 inst_7455 ( .QN(net_8940), .D(net_4741), .CK(net_16439), .RN(x6501) );
AOI22_X2 inst_8443 ( .B1(net_6601), .A1(net_6568), .A2(net_6257), .B2(net_6110), .ZN(net_3498) );
CLKBUF_X2 inst_16047 ( .A(net_15894), .Z(net_15895) );
OAI21_X2 inst_3161 ( .ZN(net_1816), .B2(net_1635), .B1(net_1264), .A(net_1108) );
CLKBUF_X2 inst_14908 ( .A(net_10052), .Z(net_14756) );
CLKBUF_X2 inst_10032 ( .A(net_9757), .Z(net_9880) );
CLKBUF_X2 inst_11462 ( .A(net_11309), .Z(net_11310) );
OR2_X4 inst_2816 ( .A1(net_5520), .ZN(net_4908), .A2(net_4898) );
XNOR2_X2 inst_276 ( .ZN(net_1032), .B(net_672), .A(net_200) );
CLKBUF_X2 inst_18640 ( .A(net_18487), .Z(net_18488) );
CLKBUF_X2 inst_13380 ( .A(net_13227), .Z(net_13228) );
NOR2_X4 inst_3339 ( .ZN(net_1483), .A1(net_1180), .A2(net_1097) );
NAND4_X2 inst_3791 ( .ZN(net_3635), .A1(net_3525), .A2(net_3524), .A3(net_3523), .A4(net_3522) );
INV_X4 inst_5297 ( .ZN(net_1598), .A(net_1597) );
XOR2_X1 inst_91 ( .A(net_7589), .Z(net_1491), .B(net_1328) );
SDFF_X2 inst_1762 ( .Q(net_7885), .D(net_7885), .SI(net_2706), .SE(net_2543), .CK(net_18034) );
SDFF_X2 inst_2023 ( .SI(net_7932), .Q(net_7932), .D(net_2717), .SE(net_2461), .CK(net_14152) );
SDFFR_X1 inst_2779 ( .D(net_7389), .Q(net_7286), .SI(net_1959), .SE(net_1327), .CK(net_15367), .RN(x6501) );
INV_X2 inst_6508 ( .A(net_7573), .ZN(net_3143) );
MUX2_X2 inst_4919 ( .S(net_8901), .A(net_8253), .Z(net_5030), .B(net_1160) );
CLKBUF_X2 inst_13250 ( .A(net_13097), .Z(net_13098) );
DFFR_X1 inst_7424 ( .QN(net_8909), .D(net_4863), .CK(net_14858), .RN(x6501) );
NAND2_X2 inst_4715 ( .ZN(net_2767), .A1(net_1787), .A2(net_1611) );
CLKBUF_X2 inst_17622 ( .A(net_17198), .Z(net_17470) );
CLKBUF_X2 inst_18625 ( .A(net_18472), .Z(net_18473) );
INV_X16 inst_6648 ( .ZN(net_6103), .A(net_3567) );
CLKBUF_X2 inst_11897 ( .A(net_11503), .Z(net_11745) );
CLKBUF_X2 inst_14079 ( .A(net_10547), .Z(net_13927) );
CLKBUF_X2 inst_16398 ( .A(net_16245), .Z(net_16246) );
AOI221_X2 inst_8851 ( .B1(net_8577), .C1(net_8466), .C2(net_6263), .B2(net_6262), .ZN(net_6223), .A(net_4254) );
AOI22_X2 inst_8075 ( .B1(net_8107), .A1(net_7767), .B2(net_6108), .A2(net_6096), .ZN(net_4069) );
CLKBUF_X2 inst_17394 ( .A(net_11164), .Z(net_17242) );
INV_X2 inst_6415 ( .ZN(net_853), .A(net_852) );
CLKBUF_X2 inst_11187 ( .A(net_11034), .Z(net_11035) );
INV_X4 inst_5161 ( .ZN(net_3178), .A(net_3158) );
CLKBUF_X2 inst_18803 ( .A(net_18650), .Z(net_18651) );
CLKBUF_X2 inst_18813 ( .A(net_18660), .Z(net_18661) );
CLKBUF_X2 inst_16754 ( .A(net_16601), .Z(net_16602) );
AOI22_X2 inst_7984 ( .B1(net_8095), .A1(net_7755), .B2(net_6108), .A2(net_6096), .ZN(net_4147) );
INV_X2 inst_6489 ( .A(net_7509), .ZN(net_556) );
XNOR2_X2 inst_266 ( .A(net_6830), .ZN(net_1112), .B(net_1029) );
SDFF_X2 inst_2051 ( .SI(net_7775), .Q(net_7775), .D(net_2655), .SE(net_2459), .CK(net_15470) );
CLKBUF_X2 inst_9288 ( .A(net_9120), .Z(net_9136) );
AOI22_X2 inst_8382 ( .B1(net_8709), .A1(net_8487), .B2(net_4350), .A2(net_4349), .ZN(net_3666) );
CLKBUF_X2 inst_18766 ( .A(net_18613), .Z(net_18614) );
CLKBUF_X2 inst_17276 ( .A(net_17123), .Z(net_17124) );
SDFF_X2 inst_1198 ( .SI(net_7300), .Q(net_7157), .D(net_7157), .SE(net_6279), .CK(net_15926) );
XNOR2_X2 inst_171 ( .B(net_2318), .ZN(net_1795), .A(net_1794) );
CLKBUF_X2 inst_17835 ( .A(net_13166), .Z(net_17683) );
CLKBUF_X2 inst_10950 ( .A(net_10797), .Z(net_10798) );
SDFF_X2 inst_374 ( .SI(net_8534), .Q(net_8534), .SE(net_3979), .D(net_3973), .CK(net_12362) );
CLKBUF_X2 inst_18023 ( .A(net_13956), .Z(net_17871) );
XOR2_X1 inst_103 ( .A(net_6835), .Z(net_1088), .B(net_990) );
CLKBUF_X2 inst_12832 ( .A(net_12679), .Z(net_12680) );
CLKBUF_X2 inst_14864 ( .A(net_14711), .Z(net_14712) );
NAND4_X2 inst_3690 ( .ZN(net_4447), .A4(net_4347), .A1(net_3827), .A2(net_3826), .A3(net_3825) );
CLKBUF_X2 inst_17372 ( .A(net_13711), .Z(net_17220) );
CLKBUF_X2 inst_10763 ( .A(net_9240), .Z(net_10611) );
INV_X2 inst_6353 ( .ZN(net_2240), .A(net_2239) );
INV_X4 inst_6061 ( .A(net_7608), .ZN(net_2493) );
CLKBUF_X2 inst_11716 ( .A(net_11563), .Z(net_11564) );
CLKBUF_X2 inst_9905 ( .A(net_9752), .Z(net_9753) );
NAND4_X2 inst_3738 ( .ZN(net_4292), .A1(net_4088), .A2(net_4087), .A3(net_4086), .A4(net_4085) );
OR2_X4 inst_2855 ( .A1(net_3187), .ZN(net_1342), .A2(net_913) );
AOI22_X2 inst_8247 ( .B1(net_8724), .A1(net_8502), .B2(net_4350), .A2(net_4349), .ZN(net_3790) );
DFF_X1 inst_6749 ( .Q(net_6758), .D(net_5618), .CK(net_10498) );
CLKBUF_X2 inst_10097 ( .A(net_9944), .Z(net_9945) );
SDFF_X2 inst_2058 ( .SI(net_7910), .Q(net_7910), .D(net_2705), .SE(net_2461), .CK(net_15800) );
SDFF_X2 inst_809 ( .SI(net_8499), .Q(net_8499), .D(net_3967), .SE(net_3884), .CK(net_13090) );
CLKBUF_X2 inst_19107 ( .A(net_18954), .Z(net_18955) );
CLKBUF_X2 inst_16609 ( .A(net_12468), .Z(net_16457) );
NAND4_X2 inst_3675 ( .A4(net_5994), .A1(net_5993), .ZN(net_4590), .A2(net_4041), .A3(net_4040) );
CLKBUF_X2 inst_15821 ( .A(net_11411), .Z(net_15669) );
AOI22_X2 inst_7816 ( .A2(net_8223), .B2(net_6144), .A1(net_4764), .ZN(net_4738), .B1(net_4666) );
SDFFR_X2 inst_2562 ( .QN(net_6352), .SE(net_2147), .D(net_2128), .SI(net_1810), .CK(net_14687), .RN(x6501) );
CLKBUF_X2 inst_14245 ( .A(net_14092), .Z(net_14093) );
SDFF_X2 inst_1022 ( .SI(net_7338), .Q(net_6679), .D(net_6679), .SE(net_3126), .CK(net_9487) );
CLKBUF_X2 inst_13925 ( .A(net_13772), .Z(net_13773) );
CLKBUF_X2 inst_15054 ( .A(net_14293), .Z(net_14902) );
CLKBUF_X2 inst_9248 ( .A(net_9066), .Z(net_9096) );
CLKBUF_X2 inst_16876 ( .A(net_9823), .Z(net_16724) );
CLKBUF_X2 inst_10416 ( .A(net_9068), .Z(net_10264) );
INV_X2 inst_6241 ( .ZN(net_4895), .A(net_4798) );
NAND3_X2 inst_3906 ( .ZN(net_5632), .A1(net_5561), .A3(net_5495), .A2(net_5370) );
AOI21_X2 inst_8928 ( .B2(net_5784), .ZN(net_5684), .A(net_5671), .B1(net_2674) );
AOI222_X1 inst_8657 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3909), .B1(net_2034), .C1(net_2033), .A1(x13863) );
CLKBUF_X2 inst_19187 ( .A(net_19034), .Z(net_19035) );
CLKBUF_X2 inst_9322 ( .A(net_9123), .Z(net_9170) );
CLKBUF_X2 inst_15103 ( .A(net_14950), .Z(net_14951) );
CLKBUF_X2 inst_10665 ( .A(net_10512), .Z(net_10513) );
CLKBUF_X2 inst_16804 ( .A(net_11673), .Z(net_16652) );
OAI22_X2 inst_2915 ( .B2(net_4221), .ZN(net_3968), .A2(net_3552), .A1(net_1464), .B1(net_668) );
CLKBUF_X2 inst_17387 ( .A(net_17234), .Z(net_17235) );
NOR3_X2 inst_3296 ( .ZN(net_1907), .A1(net_1747), .A2(net_973), .A3(net_947) );
CLKBUF_X2 inst_18129 ( .A(net_17976), .Z(net_17977) );
INV_X4 inst_6148 ( .A(net_6149), .ZN(net_6148) );
AND2_X4 inst_9135 ( .ZN(net_1415), .A2(net_802), .A1(net_183) );
CLKBUF_X2 inst_14792 ( .A(net_14639), .Z(net_14640) );
INV_X2 inst_6379 ( .A(net_1608), .ZN(net_1351) );
SDFF_X2 inst_532 ( .Q(net_8855), .D(net_8855), .SI(net_3977), .SE(net_3936), .CK(net_11095) );
OAI21_X2 inst_3164 ( .ZN(net_2703), .A(net_1661), .B1(net_1335), .B2(net_1265) );
OAI221_X2 inst_2965 ( .C2(net_3064), .B2(net_3063), .ZN(net_3062), .A(net_2880), .B1(net_2296), .C1(net_1270) );
SDFFR_X2 inst_2382 ( .SE(net_2260), .Q(net_312), .D(net_312), .CK(net_10457), .RN(x6501), .SI(x3451) );
CLKBUF_X2 inst_12228 ( .A(net_12075), .Z(net_12076) );
OAI221_X2 inst_2969 ( .C2(net_2650), .B2(net_2649), .ZN(net_2647), .A(net_2646), .C1(net_1275), .B1(net_735) );
NOR3_X2 inst_3314 ( .ZN(net_1679), .A3(net_1431), .A1(net_1148), .A2(net_859) );
CLKBUF_X2 inst_14854 ( .A(net_14701), .Z(net_14702) );
CLKBUF_X2 inst_15891 ( .A(net_15738), .Z(net_15739) );
NAND2_X4 inst_4037 ( .ZN(net_2897), .A1(net_2420), .A2(net_2331) );
CLKBUF_X2 inst_15294 ( .A(net_11800), .Z(net_15142) );
CLKBUF_X2 inst_13277 ( .A(net_13124), .Z(net_13125) );
SDFF_X2 inst_1327 ( .SI(net_7686), .Q(net_7686), .SE(net_2714), .D(net_2575), .CK(net_16005) );
CLKBUF_X2 inst_12073 ( .A(net_11263), .Z(net_11921) );
CLKBUF_X2 inst_13566 ( .A(net_13413), .Z(net_13414) );
CLKBUF_X2 inst_10598 ( .A(net_10445), .Z(net_10446) );
CLKBUF_X2 inst_11715 ( .A(net_11562), .Z(net_11563) );
CLKBUF_X2 inst_16423 ( .A(net_16270), .Z(net_16271) );
CLKBUF_X2 inst_16683 ( .A(net_15544), .Z(net_16531) );
CLKBUF_X2 inst_17969 ( .A(net_17816), .Z(net_17817) );
CLKBUF_X2 inst_16943 ( .A(net_14910), .Z(net_16791) );
INV_X4 inst_6066 ( .A(net_6311), .ZN(net_2758) );
SDFF_X2 inst_1255 ( .Q(net_8078), .D(net_8078), .SI(net_2721), .SE(net_2707), .CK(net_15782) );
CLKBUF_X2 inst_9844 ( .A(net_9691), .Z(net_9692) );
CLKBUF_X2 inst_9279 ( .A(net_9126), .Z(net_9127) );
SDFF_X2 inst_1791 ( .SI(net_8066), .Q(net_8066), .D(net_2712), .SE(net_2508), .CK(net_13747) );
NOR2_X2 inst_3420 ( .A2(net_7646), .ZN(net_3159), .A1(net_3158) );
AOI221_X2 inst_8834 ( .B1(net_8067), .C1(net_7863), .B2(net_6107), .ZN(net_6017), .C2(net_4400), .A(net_4295) );
INV_X4 inst_5064 ( .ZN(net_5919), .A(net_5872) );
CLKBUF_X2 inst_12341 ( .A(net_12188), .Z(net_12189) );
CLKBUF_X2 inst_11827 ( .A(net_10207), .Z(net_11675) );
SDFF_X2 inst_528 ( .Q(net_8884), .D(net_8884), .SI(net_3950), .SE(net_3936), .CK(net_13260) );
CLKBUF_X2 inst_9360 ( .A(net_9112), .Z(net_9208) );
CLKBUF_X2 inst_9782 ( .A(net_9629), .Z(net_9630) );
CLKBUF_X2 inst_13574 ( .A(net_13421), .Z(net_13422) );
CLKBUF_X2 inst_16244 ( .A(net_16091), .Z(net_16092) );
CLKBUF_X2 inst_17065 ( .A(net_16912), .Z(net_16913) );
CLKBUF_X2 inst_13173 ( .A(net_9388), .Z(net_13021) );
MUX2_X2 inst_4957 ( .A(net_7393), .S(net_2378), .Z(net_2366), .B(net_849) );
SDFF_X2 inst_846 ( .SI(net_8658), .Q(net_8658), .D(net_3953), .SE(net_3885), .CK(net_10227) );
CLKBUF_X2 inst_11377 ( .A(net_11224), .Z(net_11225) );
INV_X4 inst_5925 ( .A(net_8216), .ZN(net_759) );
SDFF_X2 inst_1734 ( .Q(net_7890), .D(net_7890), .SI(net_2575), .SE(net_2543), .CK(net_15962) );
DFFR_X2 inst_7036 ( .QN(net_7505), .D(net_4937), .CK(net_14511), .RN(x6501) );
CLKBUF_X2 inst_17976 ( .A(net_17823), .Z(net_17824) );
NAND2_X2 inst_4646 ( .ZN(net_2345), .A1(net_2344), .A2(net_2341) );
NOR2_X2 inst_3354 ( .ZN(net_5571), .A1(net_5412), .A2(net_5411) );
CLKBUF_X2 inst_17887 ( .A(net_17734), .Z(net_17735) );
MUX2_X2 inst_4993 ( .A(net_9026), .Z(net_3962), .B(net_3014), .S(net_622) );
CLKBUF_X2 inst_9500 ( .A(net_9347), .Z(net_9348) );
AOI22_X2 inst_8199 ( .B1(net_8755), .A1(net_8385), .A2(net_3867), .B2(net_3866), .ZN(net_3837) );
CLKBUF_X2 inst_17215 ( .A(net_17062), .Z(net_17063) );
NAND3_X2 inst_3927 ( .ZN(net_5611), .A1(net_5539), .A3(net_4648), .A2(net_4503) );
SDFFR_X1 inst_2718 ( .SI(net_9027), .Q(net_9027), .D(net_7456), .SE(net_3208), .CK(net_12933), .RN(x6501) );
XOR2_X2 inst_58 ( .B(net_6838), .A(net_990), .Z(net_964) );
NAND4_X2 inst_3633 ( .ZN(net_5335), .A2(net_4970), .A4(net_4870), .A1(net_4811), .A3(net_4580) );
CLKBUF_X2 inst_9574 ( .A(net_9128), .Z(net_9422) );
CLKBUF_X2 inst_11653 ( .A(net_11500), .Z(net_11501) );
CLKBUF_X2 inst_9775 ( .A(net_9420), .Z(net_9623) );
CLKBUF_X2 inst_13792 ( .A(net_13639), .Z(net_13640) );
SDFF_X2 inst_1469 ( .SI(net_7294), .Q(net_7151), .D(net_7151), .SE(net_6279), .CK(net_17701) );
CLKBUF_X2 inst_18806 ( .A(net_16400), .Z(net_18654) );
CLKBUF_X2 inst_10295 ( .A(net_10142), .Z(net_10143) );
CLKBUF_X2 inst_12056 ( .A(net_11903), .Z(net_11904) );
CLKBUF_X2 inst_16156 ( .A(net_16003), .Z(net_16004) );
CLKBUF_X2 inst_17949 ( .A(net_17796), .Z(net_17797) );
CLKBUF_X2 inst_12878 ( .A(net_12725), .Z(net_12726) );
CLKBUF_X2 inst_16918 ( .A(net_13859), .Z(net_16766) );
INV_X4 inst_5690 ( .ZN(net_2696), .A(net_146) );
CLKBUF_X2 inst_9592 ( .A(net_9140), .Z(net_9440) );
INV_X4 inst_5288 ( .ZN(net_1783), .A(net_1379) );
CLKBUF_X2 inst_18302 ( .A(net_12767), .Z(net_18150) );
SDFFR_X2 inst_2424 ( .D(net_2677), .SE(net_2313), .SI(net_446), .Q(net_446), .CK(net_16537), .RN(x6501) );
CLKBUF_X2 inst_15860 ( .A(net_15707), .Z(net_15708) );
NAND2_X2 inst_4517 ( .ZN(net_3875), .A2(net_3536), .A1(net_3354) );
CLKBUF_X2 inst_13719 ( .A(net_13317), .Z(net_13567) );
OAI21_X2 inst_3144 ( .ZN(net_2051), .A(net_2050), .B1(net_2049), .B2(net_2048) );
CLKBUF_X2 inst_13386 ( .A(net_9749), .Z(net_13234) );
INV_X4 inst_6124 ( .A(net_7585), .ZN(net_482) );
CLKBUF_X2 inst_11530 ( .A(net_11377), .Z(net_11378) );
NAND4_X2 inst_3666 ( .A4(net_6022), .A1(net_6021), .ZN(net_4599), .A2(net_4096), .A3(net_4095) );
SDFF_X2 inst_993 ( .D(net_7331), .SI(net_6639), .Q(net_6639), .SE(net_3123), .CK(net_11647) );
CLKBUF_X2 inst_14882 ( .A(net_14729), .Z(net_14730) );
INV_X4 inst_5177 ( .ZN(net_3153), .A(net_3022) );
INV_X2 inst_6407 ( .ZN(net_1071), .A(net_1070) );
CLKBUF_X2 inst_14590 ( .A(net_10452), .Z(net_14438) );
CLKBUF_X2 inst_17137 ( .A(net_9118), .Z(net_16985) );
CLKBUF_X2 inst_17034 ( .A(net_16881), .Z(net_16882) );
DFFR_X2 inst_7264 ( .QN(net_7358), .D(net_2006), .CK(net_11816), .RN(x6501) );
CLKBUF_X2 inst_13855 ( .A(net_13702), .Z(net_13703) );
CLKBUF_X2 inst_16646 ( .A(net_16493), .Z(net_16494) );
INV_X4 inst_5535 ( .ZN(net_822), .A(net_654) );
SDFF_X2 inst_630 ( .SI(net_8543), .Q(net_8543), .SE(net_3979), .D(net_3955), .CK(net_11006) );
INV_X4 inst_5268 ( .ZN(net_2147), .A(net_1710) );
CLKBUF_X2 inst_11796 ( .A(net_11643), .Z(net_11644) );
CLKBUF_X2 inst_9662 ( .A(net_9143), .Z(net_9510) );
SDFF_X2 inst_1273 ( .Q(net_8085), .D(net_8085), .SE(net_2707), .SI(net_2658), .CK(net_18890) );
SDFF_X2 inst_512 ( .Q(net_8865), .D(net_8865), .SI(net_3966), .SE(net_3936), .CK(net_10939) );
CLKBUF_X2 inst_11337 ( .A(net_10287), .Z(net_11185) );
CLKBUF_X2 inst_12791 ( .A(net_12638), .Z(net_12639) );
MUX2_X2 inst_4966 ( .A(net_2796), .S(net_2378), .Z(net_2357), .B(net_850) );
CLKBUF_X2 inst_14307 ( .A(net_14154), .Z(net_14155) );
CLKBUF_X2 inst_12278 ( .A(net_12125), .Z(net_12126) );
CLKBUF_X2 inst_15308 ( .A(net_9260), .Z(net_15156) );
SDFFR_X2 inst_2151 ( .Q(net_8275), .D(net_8275), .SI(net_8271), .SE(net_2996), .CK(net_18448), .RN(x6501) );
OAI21_X2 inst_3054 ( .B2(net_8235), .B1(net_4850), .ZN(net_4757), .A(net_2609) );
CLKBUF_X2 inst_15450 ( .A(net_15297), .Z(net_15298) );
CLKBUF_X2 inst_11744 ( .A(net_11591), .Z(net_11592) );
NAND2_X2 inst_4764 ( .A1(net_6340), .ZN(net_1895), .A2(net_1089) );
CLKBUF_X2 inst_18750 ( .A(net_12629), .Z(net_18598) );
CLKBUF_X2 inst_13271 ( .A(net_13118), .Z(net_13119) );
CLKBUF_X2 inst_15755 ( .A(net_12966), .Z(net_15603) );
NAND4_X2 inst_3772 ( .ZN(net_4249), .A1(net_3755), .A2(net_3754), .A3(net_3753), .A4(net_3752) );
NAND2_X2 inst_4210 ( .A1(net_7000), .ZN(net_5252), .A2(net_5249) );
SDFF_X2 inst_2043 ( .SI(net_7933), .Q(net_7933), .D(net_2711), .SE(net_2461), .CK(net_17045) );
SDFF_X2 inst_960 ( .SI(net_7318), .Q(net_6692), .D(net_6692), .SE(net_3125), .CK(net_12132) );
CLKBUF_X2 inst_16051 ( .A(net_12557), .Z(net_15899) );
SDFFR_X2 inst_2411 ( .SI(net_5946), .SE(net_2260), .Q(net_347), .D(net_347), .CK(net_9349), .RN(x6501) );
XOR2_X2 inst_38 ( .A(net_1864), .B(net_1650), .Z(net_1116) );
SDFFR_X2 inst_2601 ( .Q(net_7395), .D(net_1330), .SE(net_1136), .CK(net_18313), .RN(x6501), .SI(x4455) );
SDFF_X2 inst_381 ( .SI(net_8391), .Q(net_8391), .SE(net_3969), .D(net_3957), .CK(net_13298) );
CLKBUF_X2 inst_14846 ( .A(net_14693), .Z(net_14694) );
CLKBUF_X2 inst_9448 ( .A(net_9254), .Z(net_9296) );
NAND4_X2 inst_3837 ( .A4(net_7223), .A2(net_2767), .ZN(net_2086), .A1(net_2085), .A3(net_2084) );
DFFS_X2 inst_6876 ( .QN(net_7212), .D(net_3540), .CK(net_18927), .SN(x6501) );
DFFR_X1 inst_7577 ( .D(net_6404), .QN(net_5951), .CK(net_18008), .RN(x6501) );
CLKBUF_X2 inst_10355 ( .A(net_10202), .Z(net_10203) );
CLKBUF_X2 inst_13108 ( .A(net_9818), .Z(net_12956) );
AOI22_X2 inst_8068 ( .B1(net_7936), .A1(net_7834), .B2(net_6103), .A2(net_4398), .ZN(net_4075) );
INV_X4 inst_5496 ( .A(net_1237), .ZN(net_855) );
CLKBUF_X2 inst_18135 ( .A(net_17982), .Z(net_17983) );
INV_X4 inst_6002 ( .A(net_7640), .ZN(net_678) );
CLKBUF_X2 inst_13880 ( .A(net_13727), .Z(net_13728) );
CLKBUF_X2 inst_10228 ( .A(net_10075), .Z(net_10076) );
CLKBUF_X2 inst_14599 ( .A(net_14446), .Z(net_14447) );
CLKBUF_X2 inst_15008 ( .A(net_14855), .Z(net_14856) );
INV_X4 inst_5503 ( .A(net_1808), .ZN(net_699) );
NAND2_X2 inst_4597 ( .A1(net_6754), .A2(net_2897), .ZN(net_2844) );
SDFF_X2 inst_1188 ( .D(net_7335), .SI(net_6577), .Q(net_6577), .SE(net_3070), .CK(net_9741) );
CLKBUF_X2 inst_14579 ( .A(net_14426), .Z(net_14427) );
CLKBUF_X2 inst_13462 ( .A(net_13309), .Z(net_13310) );
CLKBUF_X2 inst_9960 ( .A(net_9756), .Z(net_9808) );
DFFS_X1 inst_6957 ( .D(net_2586), .CK(net_16577), .SN(x6501), .Q(x668) );
DFFR_X2 inst_7184 ( .QN(net_6323), .D(net_2510), .CK(net_17627), .RN(x6501) );
AOI21_X2 inst_8966 ( .A(net_7172), .ZN(net_3036), .B2(net_3035), .B1(net_1743) );
NAND3_X4 inst_3873 ( .A3(net_6185), .ZN(net_6063), .A2(net_3258), .A1(net_2328) );
AOI22_X2 inst_8363 ( .A1(net_8629), .B1(net_8444), .A2(net_3864), .B2(net_3863), .ZN(net_3685) );
CLKBUF_X2 inst_19017 ( .A(net_18864), .Z(net_18865) );
CLKBUF_X2 inst_16290 ( .A(net_15371), .Z(net_16138) );
SDFF_X2 inst_387 ( .Q(net_8818), .D(net_8818), .SI(net_3977), .SE(net_3964), .CK(net_13007) );
CLKBUF_X2 inst_18370 ( .A(net_18217), .Z(net_18218) );
NAND2_X2 inst_4601 ( .ZN(net_2888), .A2(net_2642), .A1(net_1481) );
CLKBUF_X2 inst_15416 ( .A(net_15263), .Z(net_15264) );
CLKBUF_X2 inst_14769 ( .A(net_14616), .Z(net_14617) );
CLKBUF_X2 inst_12784 ( .A(net_12631), .Z(net_12632) );
CLKBUF_X2 inst_18757 ( .A(net_9155), .Z(net_18605) );
CLKBUF_X2 inst_18711 ( .A(net_18558), .Z(net_18559) );
SDFFR_X2 inst_2129 ( .SI(net_7175), .Q(net_7175), .D(net_6426), .SE(net_4362), .CK(net_13566), .RN(x6501) );
AOI221_X2 inst_8801 ( .C2(net_6187), .B2(net_5267), .ZN(net_4835), .A(net_4834), .C1(net_191), .B1(net_171) );
INV_X4 inst_5750 ( .A(net_7242), .ZN(net_1950) );
CLKBUF_X2 inst_18714 ( .A(net_18561), .Z(net_18562) );
CLKBUF_X2 inst_11273 ( .A(net_11120), .Z(net_11121) );
CLKBUF_X2 inst_16422 ( .A(net_16269), .Z(net_16270) );
SDFF_X2 inst_1181 ( .SI(net_7323), .Q(net_6598), .D(net_6598), .SE(net_3069), .CK(net_11340) );
CLKBUF_X2 inst_18223 ( .A(net_18070), .Z(net_18071) );
AOI21_X2 inst_8986 ( .ZN(net_1884), .B2(net_1883), .B1(net_1352), .A(net_1107) );
INV_X32 inst_6165 ( .ZN(net_5443), .A(net_4904) );
INV_X8 inst_5045 ( .ZN(net_6109), .A(net_3370) );
CLKBUF_X2 inst_17863 ( .A(net_17710), .Z(net_17711) );
SDFF_X2 inst_1548 ( .Q(net_8005), .D(net_8005), .SI(net_2660), .SE(net_2542), .CK(net_14274) );
CLKBUF_X2 inst_15916 ( .A(net_15763), .Z(net_15764) );
CLKBUF_X2 inst_17100 ( .A(net_16947), .Z(net_16948) );
CLKBUF_X2 inst_9913 ( .A(net_9231), .Z(net_9761) );
CLKBUF_X2 inst_17607 ( .A(net_15364), .Z(net_17455) );
DFFR_X2 inst_7013 ( .QN(net_6304), .D(net_5720), .CK(net_14034), .RN(x6501) );
CLKBUF_X2 inst_9457 ( .A(net_9304), .Z(net_9305) );
CLKBUF_X2 inst_14255 ( .A(net_14102), .Z(net_14103) );
CLKBUF_X2 inst_10899 ( .A(net_10746), .Z(net_10747) );
INV_X4 inst_5715 ( .A(net_8916), .ZN(net_2630) );
AOI22_X2 inst_8470 ( .B1(net_6673), .A1(net_6640), .A2(net_6213), .B2(net_6138), .ZN(net_3470) );
CLKBUF_X2 inst_18338 ( .A(net_18185), .Z(net_18186) );
CLKBUF_X2 inst_10462 ( .A(net_10309), .Z(net_10310) );
AOI22_X2 inst_7799 ( .A2(net_6130), .B2(net_4965), .ZN(net_4790), .A1(net_1409), .B1(net_305) );
CLKBUF_X2 inst_16089 ( .A(net_15936), .Z(net_15937) );
CLKBUF_X2 inst_12018 ( .A(net_11865), .Z(net_11866) );
INV_X4 inst_5130 ( .ZN(net_4557), .A(net_4353) );
CLKBUF_X2 inst_14629 ( .A(net_11378), .Z(net_14477) );
CLKBUF_X2 inst_15447 ( .A(net_10389), .Z(net_15295) );
INV_X4 inst_5489 ( .ZN(net_725), .A(x3524) );
CLKBUF_X2 inst_16765 ( .A(net_16612), .Z(net_16613) );
AOI22_X2 inst_7765 ( .B1(net_6992), .A1(net_6952), .A2(net_5443), .B2(net_5442), .ZN(net_5346) );
CLKBUF_X2 inst_16453 ( .A(net_16300), .Z(net_16301) );
CLKBUF_X2 inst_14662 ( .A(net_14509), .Z(net_14510) );
AOI222_X1 inst_8682 ( .B1(net_6481), .A2(net_3296), .B2(net_3295), .C2(net_3294), .ZN(net_3290), .A1(net_3286), .C1(net_1202) );
CLKBUF_X2 inst_9760 ( .A(net_9576), .Z(net_9608) );
INV_X4 inst_5290 ( .A(net_3262), .ZN(net_1611) );
CLKBUF_X2 inst_10239 ( .A(net_10086), .Z(net_10087) );
CLKBUF_X2 inst_16468 ( .A(net_16315), .Z(net_16316) );
AOI22_X2 inst_8585 ( .B2(net_6321), .ZN(net_1792), .A2(net_1253), .B1(net_1252), .A1(x4323) );
SDFFR_X2 inst_2307 ( .SE(net_2260), .Q(net_380), .D(net_380), .CK(net_11406), .RN(x6501), .SI(x1305) );
CLKBUF_X2 inst_11611 ( .A(net_9220), .Z(net_11459) );
SDFFR_X2 inst_2611 ( .Q(net_7380), .D(net_7380), .SE(net_1136), .CK(net_18647), .RN(x6501), .SI(x4733) );
CLKBUF_X2 inst_13469 ( .A(net_11470), .Z(net_13317) );
MUX2_X2 inst_5004 ( .A(net_9037), .Z(net_3963), .B(net_3167), .S(net_622) );
CLKBUF_X2 inst_9926 ( .A(net_9773), .Z(net_9774) );
OAI21_X2 inst_2994 ( .B2(net_5902), .ZN(net_5899), .A(net_5831), .B1(net_748) );
OAI21_X2 inst_3023 ( .ZN(net_4974), .B2(net_4971), .A(net_4796), .B1(net_627) );
SDFF_X2 inst_1243 ( .Q(net_7948), .D(net_7948), .SE(net_2755), .SI(net_2708), .CK(net_15560) );
CLKBUF_X2 inst_13155 ( .A(net_13002), .Z(net_13003) );
CLKBUF_X2 inst_14970 ( .A(net_14817), .Z(net_14818) );
CLKBUF_X2 inst_9512 ( .A(net_9359), .Z(net_9360) );
CLKBUF_X2 inst_13074 ( .A(net_12921), .Z(net_12922) );
CLKBUF_X2 inst_10514 ( .A(net_10361), .Z(net_10362) );
CLKBUF_X2 inst_14639 ( .A(net_12321), .Z(net_14487) );
INV_X4 inst_5958 ( .A(net_7248), .ZN(net_1946) );
SDFF_X2 inst_1093 ( .D(net_7319), .SI(net_6495), .Q(net_6495), .SE(net_3071), .CK(net_9846) );
CLKBUF_X2 inst_14728 ( .A(net_14575), .Z(net_14576) );
NOR3_X2 inst_3271 ( .ZN(net_2416), .A1(net_2415), .A3(net_2397), .A2(net_1780) );
SDFF_X2 inst_1430 ( .SI(net_7298), .Q(net_7075), .D(net_7075), .SE(net_6280), .CK(net_18210) );
CLKBUF_X2 inst_10707 ( .A(net_10554), .Z(net_10555) );
CLKBUF_X2 inst_14516 ( .A(net_12284), .Z(net_14364) );
NOR3_X2 inst_3257 ( .ZN(net_5270), .A3(net_4973), .A1(x12843), .A2(x12810) );
CLKBUF_X2 inst_10759 ( .A(net_9275), .Z(net_10607) );
CLKBUF_X2 inst_14081 ( .A(net_13928), .Z(net_13929) );
CLKBUF_X2 inst_11498 ( .A(net_11321), .Z(net_11346) );
CLKBUF_X2 inst_16543 ( .A(net_16390), .Z(net_16391) );
CLKBUF_X2 inst_9979 ( .A(net_9691), .Z(net_9827) );
SDFF_X2 inst_763 ( .Q(net_8806), .D(net_8806), .SI(net_3953), .SE(net_3879), .CK(net_10240) );
SDFFR_X2 inst_2330 ( .SI(net_7367), .D(net_2741), .SE(net_2740), .QN(net_278), .CK(net_16419), .RN(x6501) );
DFFR_X1 inst_7377 ( .QN(net_6316), .D(net_5915), .CK(net_16952), .RN(x6501) );
NAND4_X2 inst_3636 ( .ZN(net_5276), .A4(net_4867), .A2(net_4673), .A1(net_4538), .A3(net_4488) );
CLKBUF_X2 inst_11069 ( .A(net_9467), .Z(net_10917) );
CLKBUF_X2 inst_14018 ( .A(net_13865), .Z(net_13866) );
CLKBUF_X2 inst_13754 ( .A(net_13601), .Z(net_13602) );
CLKBUF_X2 inst_15970 ( .A(net_15817), .Z(net_15818) );
CLKBUF_X2 inst_17185 ( .A(net_12052), .Z(net_17033) );
SDFF_X2 inst_537 ( .Q(net_8678), .D(net_8678), .SI(net_3962), .SE(net_3935), .CK(net_12992) );
INV_X4 inst_5069 ( .ZN(net_5859), .A(net_5813) );
CLKBUF_X2 inst_17935 ( .A(net_17782), .Z(net_17783) );
DFFR_X2 inst_7141 ( .QN(net_7343), .D(net_2962), .CK(net_11617), .RN(x6501) );
CLKBUF_X2 inst_14977 ( .A(net_14824), .Z(net_14825) );
CLKBUF_X2 inst_15232 ( .A(net_15079), .Z(net_15080) );
CLKBUF_X2 inst_14341 ( .A(net_13323), .Z(net_14189) );
AOI22_X2 inst_8431 ( .B1(net_6598), .A1(net_6565), .A2(net_6257), .B2(net_6110), .ZN(net_3510) );
CLKBUF_X2 inst_10786 ( .A(net_10633), .Z(net_10634) );
NAND3_X2 inst_3950 ( .ZN(net_4273), .A3(net_4216), .A2(net_3928), .A1(net_3927) );
AOI221_X2 inst_8863 ( .ZN(net_2102), .A(net_1628), .B1(net_1527), .C2(net_1526), .C1(net_1337), .B2(net_1263) );
NAND2_X2 inst_4288 ( .A1(net_7009), .A2(net_5249), .ZN(net_5172) );
SDFF_X2 inst_869 ( .Q(net_8579), .D(net_8579), .SI(net_3942), .SE(net_3878), .CK(net_12782) );
CLKBUF_X2 inst_10671 ( .A(net_10518), .Z(net_10519) );
SDFFR_X1 inst_2646 ( .D(net_6769), .SE(net_4506), .CK(net_9247), .RN(x6501), .SI(x1804), .Q(x1804) );
CLKBUF_X2 inst_18321 ( .A(net_9484), .Z(net_18169) );
INV_X2 inst_6543 ( .A(net_7622), .ZN(net_1315) );
CLKBUF_X2 inst_18493 ( .A(net_18340), .Z(net_18341) );
CLKBUF_X2 inst_17824 ( .A(net_17671), .Z(net_17672) );
CLKBUF_X2 inst_13229 ( .A(net_13076), .Z(net_13077) );
CLKBUF_X2 inst_9753 ( .A(net_9600), .Z(net_9601) );
CLKBUF_X2 inst_13649 ( .A(net_13496), .Z(net_13497) );
NOR3_X2 inst_3267 ( .A3(net_2963), .ZN(net_2783), .A2(net_2290), .A1(net_1915) );
CLKBUF_X2 inst_9849 ( .A(net_9696), .Z(net_9697) );
OAI211_X2 inst_3205 ( .C2(net_5036), .ZN(net_2635), .B(net_2154), .A(net_1516), .C1(net_1174) );
CLKBUF_X2 inst_14315 ( .A(net_11759), .Z(net_14163) );
CLKBUF_X2 inst_17109 ( .A(net_16956), .Z(net_16957) );
INV_X4 inst_6048 ( .A(net_7645), .ZN(net_1637) );
AOI21_X2 inst_8945 ( .B2(net_5871), .ZN(net_5603), .A(net_5602), .B1(x563) );
SDFF_X2 inst_612 ( .SI(net_8374), .Q(net_8374), .D(net_3977), .SE(net_3969), .CK(net_10764) );
CLKBUF_X2 inst_12505 ( .A(net_12352), .Z(net_12353) );
INV_X2 inst_6185 ( .ZN(net_5834), .A(net_5780) );
SDFF_X2 inst_1692 ( .Q(net_8023), .D(net_8023), .SI(net_2720), .SE(net_2545), .CK(net_15261) );
CLKBUF_X2 inst_15875 ( .A(net_13276), .Z(net_15723) );
NAND3_X2 inst_3986 ( .ZN(net_1913), .A3(net_1543), .A1(net_1203), .A2(net_981) );
CLKBUF_X2 inst_13137 ( .A(net_12984), .Z(net_12985) );
DFFR_X2 inst_7275 ( .QN(net_7306), .D(net_1875), .CK(net_18338), .RN(x6501) );
CLKBUF_X2 inst_14328 ( .A(net_14175), .Z(net_14176) );
CLKBUF_X2 inst_10819 ( .A(net_10666), .Z(net_10667) );
CLKBUF_X2 inst_14535 ( .A(net_14382), .Z(net_14383) );
SDFFR_X2 inst_2455 ( .D(net_2666), .SE(net_2313), .SI(net_439), .Q(net_439), .CK(net_16412), .RN(x6501) );
CLKBUF_X2 inst_18157 ( .A(net_18004), .Z(net_18005) );
CLKBUF_X2 inst_12923 ( .A(net_12770), .Z(net_12771) );
CLKBUF_X2 inst_10575 ( .A(net_10422), .Z(net_10423) );
CLKBUF_X2 inst_15690 ( .A(net_12881), .Z(net_15538) );
CLKBUF_X2 inst_17570 ( .A(net_17417), .Z(net_17418) );
DFF_X1 inst_6724 ( .Q(net_6770), .D(net_5645), .CK(net_9262) );
CLKBUF_X2 inst_11581 ( .A(net_11417), .Z(net_11429) );
NAND2_X2 inst_4828 ( .ZN(net_1331), .A2(net_1101), .A1(net_713) );
CLKBUF_X2 inst_18258 ( .A(net_18105), .Z(net_18106) );
INV_X4 inst_5218 ( .A(net_5044), .ZN(net_4803) );
INV_X4 inst_5389 ( .ZN(net_2760), .A(net_1090) );
CLKBUF_X2 inst_17152 ( .A(net_16999), .Z(net_17000) );
SDFF_X2 inst_885 ( .Q(net_8589), .D(net_8589), .SI(net_3976), .SE(net_3878), .CK(net_12778) );
CLKBUF_X2 inst_15995 ( .A(net_15842), .Z(net_15843) );
CLKBUF_X2 inst_18509 ( .A(net_18356), .Z(net_18357) );
CLKBUF_X2 inst_17796 ( .A(net_17643), .Z(net_17644) );
INV_X4 inst_5803 ( .A(net_7602), .ZN(net_1340) );
CLKBUF_X2 inst_10748 ( .A(net_10595), .Z(net_10596) );
CLKBUF_X2 inst_18314 ( .A(net_18161), .Z(net_18162) );
NOR2_X2 inst_3610 ( .A2(net_8965), .A1(net_8964), .ZN(net_1588) );
OAI21_X2 inst_2999 ( .B2(net_5902), .ZN(net_5894), .A(net_5826), .B1(net_684) );
CLKBUF_X2 inst_13097 ( .A(net_12944), .Z(net_12945) );
AOI22_X2 inst_8351 ( .B1(net_8775), .A1(net_8405), .A2(net_3867), .B2(net_3866), .ZN(net_3697) );
CLKBUF_X2 inst_12822 ( .A(net_12669), .Z(net_12670) );
AOI22_X2 inst_8188 ( .B1(net_8791), .A1(net_8532), .ZN(net_6242), .A2(net_3861), .B2(net_3860) );
INV_X4 inst_5956 ( .A(net_5954), .ZN(net_767) );
CLKBUF_X2 inst_17750 ( .A(net_14693), .Z(net_17598) );
INV_X4 inst_5305 ( .ZN(net_1498), .A(net_1367) );
NAND2_X2 inst_4156 ( .ZN(net_5359), .A2(net_5206), .A1(net_5099) );
CLKBUF_X2 inst_9875 ( .A(net_9722), .Z(net_9723) );
CLKBUF_X2 inst_16896 ( .A(net_16743), .Z(net_16744) );
XNOR2_X2 inst_200 ( .ZN(net_1544), .B(net_1204), .A(net_1191) );
CLKBUF_X2 inst_11986 ( .A(net_9443), .Z(net_11834) );
CLKBUF_X2 inst_16490 ( .A(net_16156), .Z(net_16338) );
CLKBUF_X2 inst_17649 ( .A(net_17496), .Z(net_17497) );
NAND2_X2 inst_4373 ( .A1(net_7074), .A2(net_5162), .ZN(net_5084) );
AND2_X2 inst_9198 ( .ZN(net_1580), .A1(net_1340), .A2(net_1339) );
CLKBUF_X2 inst_9939 ( .A(net_9093), .Z(net_9787) );
CLKBUF_X2 inst_18463 ( .A(net_18310), .Z(net_18311) );
CLKBUF_X2 inst_16094 ( .A(net_15941), .Z(net_15942) );
CLKBUF_X2 inst_18434 ( .A(net_18281), .Z(net_18282) );
SDFF_X2 inst_1750 ( .Q(net_7894), .D(net_7894), .SI(net_2718), .SE(net_2543), .CK(net_18762) );
INV_X4 inst_5242 ( .A(net_2159), .ZN(net_1965) );
CLKBUF_X2 inst_10155 ( .A(net_10002), .Z(net_10003) );
AOI22_X2 inst_7758 ( .B1(net_6986), .A1(net_6946), .A2(net_5443), .B2(net_5442), .ZN(net_5374) );
CLKBUF_X2 inst_16185 ( .A(net_16032), .Z(net_16033) );
CLKBUF_X2 inst_9569 ( .A(net_9308), .Z(net_9417) );
CLKBUF_X2 inst_17528 ( .A(net_17375), .Z(net_17376) );
CLKBUF_X2 inst_12294 ( .A(net_12141), .Z(net_12142) );
NOR2_X2 inst_3499 ( .ZN(net_1896), .A1(net_1895), .A2(net_1894) );
SDFF_X2 inst_893 ( .Q(net_8567), .D(net_8567), .SI(net_3962), .SE(net_3878), .CK(net_10131) );
AOI22_X2 inst_8128 ( .A1(net_7947), .B1(net_7777), .A2(net_6092), .B2(net_6091), .ZN(net_4021) );
CLKBUF_X2 inst_15711 ( .A(net_15558), .Z(net_15559) );
CLKBUF_X2 inst_15435 ( .A(net_15282), .Z(net_15283) );
CLKBUF_X2 inst_17923 ( .A(net_14458), .Z(net_17771) );
SDFF_X2 inst_569 ( .Q(net_8833), .D(net_8833), .SE(net_3964), .SI(net_3958), .CK(net_12272) );
AND2_X2 inst_9209 ( .A2(net_1489), .A1(net_970), .ZN(net_837) );
CLKBUF_X2 inst_12763 ( .A(net_9633), .Z(net_12611) );
CLKBUF_X2 inst_14730 ( .A(net_14577), .Z(net_14578) );
CLKBUF_X2 inst_15440 ( .A(net_15287), .Z(net_15288) );
CLKBUF_X2 inst_14451 ( .A(net_14298), .Z(net_14299) );
CLKBUF_X2 inst_12554 ( .A(net_12401), .Z(net_12402) );
CLKBUF_X2 inst_16328 ( .A(net_16175), .Z(net_16176) );
CLKBUF_X2 inst_18555 ( .A(net_15688), .Z(net_18403) );
NAND2_X2 inst_4220 ( .A1(net_7014), .A2(net_5249), .ZN(net_5240) );
SDFF_X2 inst_522 ( .Q(net_8877), .D(net_8877), .SI(net_3954), .SE(net_3936), .CK(net_10073) );
CLKBUF_X2 inst_18658 ( .A(net_18505), .Z(net_18506) );
INV_X8 inst_5040 ( .ZN(net_6097), .A(net_3565) );
CLKBUF_X2 inst_19172 ( .A(net_19019), .Z(net_19020) );
AND4_X2 inst_9037 ( .A1(net_2315), .ZN(net_2182), .A3(net_2181), .A4(net_2046), .A2(net_1865) );
CLKBUF_X2 inst_12408 ( .A(net_12255), .Z(net_12256) );
CLKBUF_X2 inst_14458 ( .A(net_14305), .Z(net_14306) );
CLKBUF_X2 inst_9842 ( .A(net_9689), .Z(net_9690) );
OR3_X2 inst_2809 ( .A2(net_6322), .A1(net_4924), .A3(net_2767), .ZN(net_2080) );
CLKBUF_X2 inst_9654 ( .A(net_9501), .Z(net_9502) );
CLKBUF_X2 inst_14011 ( .A(net_13858), .Z(net_13859) );
CLKBUF_X2 inst_15147 ( .A(net_14994), .Z(net_14995) );
CLKBUF_X2 inst_12478 ( .A(net_12325), .Z(net_12326) );
CLKBUF_X2 inst_17076 ( .A(net_16923), .Z(net_16924) );
CLKBUF_X2 inst_13141 ( .A(net_10203), .Z(net_12989) );
CLKBUF_X2 inst_12797 ( .A(net_12644), .Z(net_12645) );
CLKBUF_X2 inst_18273 ( .A(net_16332), .Z(net_18121) );
DFFS_X1 inst_6936 ( .D(net_6145), .CK(net_13654), .SN(x6501), .Q(x703) );
CLKBUF_X2 inst_18401 ( .A(net_18248), .Z(net_18249) );
CLKBUF_X2 inst_17497 ( .A(net_17344), .Z(net_17345) );
DFFS_X1 inst_6911 ( .D(net_5885), .CK(net_13818), .SN(x6501), .Q(x20) );
AND2_X4 inst_9144 ( .A2(net_7403), .A1(net_7399), .ZN(net_1504) );
CLKBUF_X2 inst_18662 ( .A(net_17534), .Z(net_18510) );
CLKBUF_X2 inst_11131 ( .A(net_10978), .Z(net_10979) );
AOI21_X2 inst_8997 ( .B1(net_7626), .B2(net_7625), .ZN(net_2959), .A(net_1315) );
INV_X2 inst_6493 ( .ZN(net_552), .A(x13193) );
CLKBUF_X2 inst_14779 ( .A(net_12084), .Z(net_14627) );
CLKBUF_X2 inst_16603 ( .A(net_15766), .Z(net_16451) );
SDFF_X2 inst_719 ( .SI(net_8640), .Q(net_8640), .D(net_3960), .SE(net_3885), .CK(net_11062) );
CLKBUF_X2 inst_15699 ( .A(net_15546), .Z(net_15547) );
CLKBUF_X2 inst_10195 ( .A(net_9403), .Z(net_10043) );
NAND2_X2 inst_4166 ( .ZN(net_5345), .A1(net_5199), .A2(net_4992) );
CLKBUF_X2 inst_18182 ( .A(net_14303), .Z(net_18030) );
CLKBUF_X2 inst_18234 ( .A(net_14194), .Z(net_18082) );
NAND3_X4 inst_3868 ( .A1(net_6260), .A3(net_6190), .A2(net_4816), .ZN(net_4815) );
AOI222_X1 inst_8695 ( .C2(net_4889), .B2(net_4888), .A1(net_4803), .ZN(net_3204), .C1(net_3203), .B1(net_3137), .A2(net_3013) );
CLKBUF_X2 inst_17574 ( .A(net_14000), .Z(net_17422) );
SDFF_X2 inst_1134 ( .D(net_7341), .SI(net_6583), .Q(net_6583), .SE(net_3070), .CK(net_11868) );
NOR2_X2 inst_3546 ( .A1(net_7490), .ZN(net_1677), .A2(net_1320) );
INV_X4 inst_5748 ( .ZN(net_2965), .A(net_289) );
SDFF_X2 inst_1144 ( .SI(net_7324), .Q(net_6599), .D(net_6599), .SE(net_3069), .CK(net_12073) );
INV_X4 inst_5165 ( .ZN(net_3158), .A(net_3081) );
INV_X2 inst_6426 ( .A(net_1271), .ZN(net_736) );
INV_X4 inst_5366 ( .A(net_2408), .ZN(net_1137) );
INV_X4 inst_5551 ( .A(net_1886), .ZN(net_878) );
CLKBUF_X2 inst_17599 ( .A(net_17446), .Z(net_17447) );
SDFFR_X2 inst_2568 ( .Q(net_6384), .D(net_6384), .SE(net_2147), .SI(net_2073), .CK(net_18229), .RN(x6501) );
SDFFR_X2 inst_2295 ( .D(net_2758), .SE(net_2757), .SI(net_470), .Q(net_470), .CK(net_13958), .RN(x6501) );
CLKBUF_X2 inst_17168 ( .A(net_12576), .Z(net_17016) );
CLKBUF_X2 inst_13021 ( .A(net_12868), .Z(net_12869) );
CLKBUF_X2 inst_17759 ( .A(net_17606), .Z(net_17607) );
CLKBUF_X2 inst_19039 ( .A(net_18886), .Z(net_18887) );
NOR2_X2 inst_3532 ( .ZN(net_1629), .A1(net_1365), .A2(net_992) );
OAI21_X2 inst_3028 ( .B2(net_4971), .ZN(net_4939), .A(net_4839), .B1(net_715) );
AND2_X2 inst_9190 ( .A2(net_2181), .ZN(net_2081), .A1(net_1104) );
NAND4_X2 inst_3854 ( .ZN(net_1557), .A3(net_1096), .A2(net_1047), .A4(net_997), .A1(net_961) );
CLKBUF_X2 inst_9432 ( .A(net_9213), .Z(net_9280) );
CLKBUF_X2 inst_10881 ( .A(net_10728), .Z(net_10729) );
DFFR_X2 inst_7089 ( .QN(net_7214), .D(net_3539), .CK(net_18964), .RN(x6501) );
SDFF_X2 inst_1530 ( .Q(net_7907), .D(net_7907), .SI(net_2703), .SE(net_2543), .CK(net_14010) );
CLKBUF_X2 inst_18004 ( .A(net_17851), .Z(net_17852) );
INV_X4 inst_5421 ( .ZN(net_4671), .A(net_857) );
CLKBUF_X2 inst_17091 ( .A(net_16938), .Z(net_16939) );
INV_X2 inst_6308 ( .ZN(net_3896), .A(net_3593) );
CLKBUF_X2 inst_11599 ( .A(net_11446), .Z(net_11447) );
CLKBUF_X2 inst_18816 ( .A(net_12642), .Z(net_18664) );
INV_X4 inst_5948 ( .A(net_8912), .ZN(net_4669) );
CLKBUF_X2 inst_9340 ( .A(net_9187), .Z(net_9188) );
INV_X2 inst_6282 ( .ZN(net_4219), .A(net_3932) );
CLKBUF_X2 inst_10076 ( .A(net_9923), .Z(net_9924) );
CLKBUF_X2 inst_10955 ( .A(net_10802), .Z(net_10803) );
CLKBUF_X2 inst_13318 ( .A(net_9461), .Z(net_13166) );
CLKBUF_X2 inst_12111 ( .A(net_9285), .Z(net_11959) );
CLKBUF_X2 inst_17598 ( .A(net_12846), .Z(net_17446) );
CLKBUF_X2 inst_19026 ( .A(net_12953), .Z(net_18874) );
CLKBUF_X2 inst_13876 ( .A(net_13723), .Z(net_13724) );
CLKBUF_X2 inst_18477 ( .A(net_18324), .Z(net_18325) );
CLKBUF_X2 inst_17051 ( .A(net_16898), .Z(net_16899) );
CLKBUF_X2 inst_12586 ( .A(net_9069), .Z(net_12434) );
INV_X2 inst_6244 ( .ZN(net_4862), .A(net_4765) );
AOI221_X2 inst_8753 ( .C2(net_6455), .C1(net_5654), .B2(net_5595), .ZN(net_5593), .A(net_5327), .B1(net_337) );
NAND2_X2 inst_4174 ( .ZN(net_5334), .A2(net_5194), .A1(net_5081) );
CLKBUF_X2 inst_17841 ( .A(net_14460), .Z(net_17689) );
CLKBUF_X2 inst_15133 ( .A(net_14980), .Z(net_14981) );
INV_X2 inst_6369 ( .ZN(net_4389), .A(net_1713) );
SDFFR_X2 inst_2502 ( .Q(net_9002), .D(net_9002), .SI(net_2628), .SE(net_2562), .CK(net_13672), .RN(x6501) );
CLKBUF_X2 inst_17473 ( .A(net_17320), .Z(net_17321) );
AND2_X4 inst_9114 ( .ZN(net_1902), .A2(net_1732), .A1(net_1513) );
CLKBUF_X2 inst_11233 ( .A(net_9133), .Z(net_11081) );
NAND3_X2 inst_3974 ( .A3(net_5582), .A2(net_3162), .ZN(net_2252), .A1(net_1999) );
CLKBUF_X2 inst_17425 ( .A(net_17272), .Z(net_17273) );
CLKBUF_X2 inst_13290 ( .A(net_13137), .Z(net_13138) );
CLKBUF_X2 inst_12601 ( .A(net_11663), .Z(net_12449) );
XNOR2_X2 inst_213 ( .ZN(net_1448), .B(net_1340), .A(net_1339) );
CLKBUF_X2 inst_11501 ( .A(net_11348), .Z(net_11349) );
CLKBUF_X2 inst_18167 ( .A(net_18014), .Z(net_18015) );
CLKBUF_X2 inst_18408 ( .A(net_18255), .Z(net_18256) );
XNOR2_X2 inst_205 ( .ZN(net_1538), .B(net_944), .A(net_928) );
SDFF_X2 inst_1645 ( .SI(net_7723), .Q(net_7723), .D(net_2722), .SE(net_2559), .CK(net_15984) );
AOI22_X2 inst_7904 ( .A2(net_5538), .ZN(net_4523), .B1(net_4522), .B2(net_4388), .A1(net_419) );
NAND4_X2 inst_3722 ( .ZN(net_4308), .A1(net_4184), .A2(net_4183), .A3(net_4182), .A4(net_4181) );
AOI22_X2 inst_8043 ( .B1(net_8171), .A1(net_7729), .B2(net_6101), .A2(net_6095), .ZN(net_6022) );
INV_X4 inst_5410 ( .ZN(net_2033), .A(net_874) );
NAND2_X2 inst_4311 ( .A1(net_7136), .A2(net_5166), .ZN(net_5146) );
CLKBUF_X2 inst_15618 ( .A(net_15465), .Z(net_15466) );
CLKBUF_X2 inst_14469 ( .A(net_14316), .Z(net_14317) );
CLKBUF_X2 inst_14916 ( .A(net_12479), .Z(net_14764) );
INV_X4 inst_5173 ( .ZN(net_2966), .A(net_2914) );
CLKBUF_X2 inst_14117 ( .A(net_12015), .Z(net_13965) );
CLKBUF_X2 inst_15388 ( .A(net_15235), .Z(net_15236) );
INV_X2 inst_6464 ( .A(net_8899), .ZN(net_2205) );
OAI221_X2 inst_2951 ( .ZN(net_4955), .B1(net_4954), .B2(net_4849), .A(net_4664), .C2(net_4559), .C1(net_817) );
AND2_X2 inst_9176 ( .A2(net_6188), .ZN(net_2390), .A1(x3327) );
NAND3_X2 inst_3890 ( .ZN(net_5648), .A1(net_5577), .A3(net_5511), .A2(net_5434) );
CLKBUF_X2 inst_13526 ( .A(net_13373), .Z(net_13374) );
CLKBUF_X2 inst_10209 ( .A(net_10056), .Z(net_10057) );
SDFFR_X2 inst_2535 ( .SI(net_7260), .Q(net_7260), .D(net_2129), .SE(net_1379), .CK(net_15033), .RN(x6501) );
NAND2_X2 inst_4569 ( .ZN(net_3122), .A1(net_3068), .A2(net_3031) );
CLKBUF_X2 inst_18873 ( .A(net_18720), .Z(net_18721) );
CLKBUF_X2 inst_12393 ( .A(net_12240), .Z(net_12241) );
NAND2_X2 inst_4480 ( .A2(net_4881), .ZN(net_4498), .A1(net_244) );
HA_X1 inst_6676 ( .A(net_3309), .S(net_3106), .CO(net_3105), .B(net_2926) );
CLKBUF_X2 inst_10723 ( .A(net_10570), .Z(net_10571) );
CLKBUF_X2 inst_9378 ( .A(net_9225), .Z(net_9226) );
CLKBUF_X2 inst_18058 ( .A(net_17905), .Z(net_17906) );
CLKBUF_X2 inst_17536 ( .A(net_15785), .Z(net_17384) );
INV_X4 inst_5639 ( .A(net_7412), .ZN(net_1457) );
NOR2_X2 inst_3502 ( .A2(net_2318), .ZN(net_2279), .A1(net_1862) );
NOR2_X2 inst_3473 ( .ZN(net_5028), .A2(net_5027), .A1(net_1349) );
CLKBUF_X2 inst_14584 ( .A(net_10663), .Z(net_14432) );
CLKBUF_X2 inst_18160 ( .A(net_18007), .Z(net_18008) );
INV_X4 inst_6018 ( .ZN(net_509), .A(net_157) );
CLKBUF_X2 inst_9942 ( .A(net_9773), .Z(net_9790) );
CLKBUF_X2 inst_14644 ( .A(net_12617), .Z(net_14492) );
AOI22_X2 inst_8502 ( .B1(net_6681), .A1(net_6648), .A2(net_6213), .B2(net_6138), .ZN(net_3438) );
CLKBUF_X2 inst_17556 ( .A(net_17403), .Z(net_17404) );
INV_X4 inst_5822 ( .A(net_5961), .ZN(x2908) );
CLKBUF_X2 inst_19123 ( .A(net_18970), .Z(net_18971) );
INV_X2 inst_6448 ( .A(net_6359), .ZN(net_2136) );
CLKBUF_X2 inst_16013 ( .A(net_15860), .Z(net_15861) );
SDFF_X2 inst_348 ( .Q(net_8744), .D(net_8744), .SE(net_3982), .SI(net_3977), .CK(net_10779) );
AOI221_X4 inst_8737 ( .B1(net_8820), .C1(net_8339), .C2(net_6265), .B2(net_6253), .ZN(net_4329), .A(net_4235) );
INV_X4 inst_5123 ( .A(net_4624), .ZN(net_4417) );
SDFFR_X1 inst_2686 ( .SI(net_7548), .SE(net_5043), .CK(net_12756), .RN(x6501), .Q(x3954), .D(x3954) );
CLKBUF_X2 inst_14911 ( .A(net_14758), .Z(net_14759) );
CLKBUF_X2 inst_10774 ( .A(net_9644), .Z(net_10622) );
NAND4_X2 inst_3740 ( .ZN(net_4290), .A1(net_4076), .A2(net_4075), .A3(net_4074), .A4(net_4073) );
SDFFR_X2 inst_2293 ( .SI(net_7378), .SE(net_2793), .Q(net_237), .D(net_237), .CK(net_17822), .RN(x6501) );
CLKBUF_X2 inst_9600 ( .A(net_9447), .Z(net_9448) );
CLKBUF_X2 inst_11299 ( .A(net_11146), .Z(net_11147) );
CLKBUF_X2 inst_18108 ( .A(net_17955), .Z(net_17956) );
SDFF_X2 inst_645 ( .SI(net_8528), .Q(net_8528), .SE(net_3979), .D(net_3946), .CK(net_11076) );
CLKBUF_X2 inst_13299 ( .A(net_13146), .Z(net_13147) );
CLKBUF_X2 inst_15615 ( .A(net_15462), .Z(net_15463) );
OAI21_X2 inst_3041 ( .B2(net_8232), .B1(net_4928), .ZN(net_4820), .A(net_3053) );
CLKBUF_X2 inst_14967 ( .A(net_14814), .Z(net_14815) );
SDFFR_X1 inst_2719 ( .SI(net_9028), .Q(net_9028), .D(net_7457), .SE(net_3208), .CK(net_10677), .RN(x6501) );
SDFFR_X2 inst_2352 ( .D(net_2729), .SE(net_2313), .SI(net_469), .Q(net_469), .CK(net_13952), .RN(x6501) );
XNOR2_X2 inst_269 ( .A(net_8255), .B(net_1206), .ZN(net_1051) );
DFFS_X2 inst_6864 ( .QN(net_8970), .D(net_5282), .CK(net_17622), .SN(x6501) );
CLKBUF_X2 inst_17125 ( .A(net_16972), .Z(net_16973) );
CLKBUF_X2 inst_12534 ( .A(net_12381), .Z(net_12382) );
CLKBUF_X2 inst_14278 ( .A(net_14125), .Z(net_14126) );
CLKBUF_X2 inst_18383 ( .A(net_18230), .Z(net_18231) );
CLKBUF_X2 inst_15947 ( .A(net_15794), .Z(net_15795) );
CLKBUF_X2 inst_9796 ( .A(net_9643), .Z(net_9644) );
SDFF_X2 inst_514 ( .Q(net_8867), .D(net_8867), .SI(net_3973), .SE(net_3936), .CK(net_12345) );
SDFF_X2 inst_1541 ( .Q(net_7977), .D(net_7977), .SI(net_2585), .SE(net_2542), .CK(net_15836) );
CLKBUF_X2 inst_12707 ( .A(net_12554), .Z(net_12555) );
CLKBUF_X2 inst_15867 ( .A(net_14504), .Z(net_15715) );
NAND2_X2 inst_4236 ( .A1(net_7021), .A2(net_5249), .ZN(net_5224) );
CLKBUF_X2 inst_16828 ( .A(net_16675), .Z(net_16676) );
CLKBUF_X2 inst_12952 ( .A(net_10612), .Z(net_12800) );
CLKBUF_X2 inst_14061 ( .A(net_13908), .Z(net_13909) );
NAND2_X2 inst_4656 ( .A1(net_2641), .A2(net_2334), .ZN(net_2272) );
CLKBUF_X2 inst_10658 ( .A(net_10505), .Z(net_10506) );
CLKBUF_X2 inst_14358 ( .A(net_14205), .Z(net_14206) );
INV_X4 inst_5621 ( .A(net_8924), .ZN(net_2592) );
CLKBUF_X2 inst_10636 ( .A(net_10158), .Z(net_10484) );
CLKBUF_X2 inst_11585 ( .A(net_11432), .Z(net_11433) );
NOR2_X2 inst_3432 ( .A2(net_3093), .ZN(net_3077), .A1(net_1448) );
CLKBUF_X2 inst_14047 ( .A(net_9397), .Z(net_13895) );
CLKBUF_X2 inst_15760 ( .A(net_15607), .Z(net_15608) );
CLKBUF_X2 inst_13984 ( .A(net_13831), .Z(net_13832) );
CLKBUF_X2 inst_15211 ( .A(net_13071), .Z(net_15059) );
AOI21_X2 inst_8959 ( .ZN(net_4957), .B1(net_4926), .A(net_4638), .B2(net_1990) );
DFFS_X2 inst_6881 ( .Q(net_8255), .D(net_3221), .CK(net_18479), .SN(x6501) );
NAND4_X2 inst_3840 ( .ZN(net_2224), .A2(net_2181), .A1(net_1870), .A3(net_1772), .A4(net_1703) );
AOI21_X2 inst_8905 ( .B2(net_5871), .ZN(net_5759), .A(net_5758), .B1(net_2726) );
CLKBUF_X2 inst_9477 ( .A(net_9324), .Z(net_9325) );
CLKBUF_X2 inst_13852 ( .A(net_13699), .Z(net_13700) );
CLKBUF_X2 inst_16695 ( .A(net_9847), .Z(net_16543) );
DFFR_X2 inst_6973 ( .QN(net_5969), .D(net_5913), .CK(net_11564), .RN(x6501) );
INV_X4 inst_5333 ( .ZN(net_1461), .A(net_1343) );
CLKBUF_X2 inst_17553 ( .A(net_17400), .Z(net_17401) );
DFFR_X2 inst_7170 ( .D(net_2578), .QN(net_341), .CK(net_11614), .RN(x6501) );
MUX2_X2 inst_4944 ( .B(net_7481), .A(net_2760), .Z(net_2524), .S(net_2343) );
CLKBUF_X2 inst_13971 ( .A(net_12250), .Z(net_13819) );
CLKBUF_X2 inst_10975 ( .A(net_9387), .Z(net_10823) );
CLKBUF_X2 inst_10259 ( .A(net_10106), .Z(net_10107) );
XNOR2_X2 inst_312 ( .ZN(net_957), .A(net_956), .B(net_955) );
CLKBUF_X2 inst_13429 ( .A(net_13276), .Z(net_13277) );
CLKBUF_X2 inst_9554 ( .A(net_9122), .Z(net_9402) );
CLKBUF_X2 inst_17829 ( .A(net_17676), .Z(net_17677) );
XNOR2_X2 inst_309 ( .A(net_4621), .ZN(net_962), .B(net_487) );
NOR2_X2 inst_3416 ( .A2(net_6080), .ZN(net_3367), .A1(net_3179) );
CLKBUF_X2 inst_13765 ( .A(net_13612), .Z(net_13613) );
CLKBUF_X2 inst_9365 ( .A(net_9212), .Z(net_9213) );
DFFR_X2 inst_7265 ( .QN(net_7210), .D(net_2026), .CK(net_18946), .RN(x6501) );
AOI22_X2 inst_8038 ( .B1(net_8102), .A1(net_7762), .B2(net_6108), .A2(net_6096), .ZN(net_4101) );
SDFFR_X1 inst_2694 ( .SI(net_7556), .SE(net_5043), .CK(net_12732), .RN(x6501), .Q(x3830), .D(x3830) );
CLKBUF_X2 inst_9833 ( .A(net_9680), .Z(net_9681) );
CLKBUF_X2 inst_15207 ( .A(net_15019), .Z(net_15055) );
SDFF_X2 inst_1968 ( .D(net_7293), .SI(net_6990), .Q(net_6990), .SE(net_6283), .CK(net_17659) );
CLKBUF_X2 inst_12983 ( .A(net_9747), .Z(net_12831) );
CLKBUF_X2 inst_12168 ( .A(net_12015), .Z(net_12016) );
SDFF_X2 inst_1330 ( .SI(net_7688), .Q(net_7688), .SE(net_2714), .D(net_2590), .CK(net_15624) );
CLKBUF_X2 inst_12038 ( .A(net_11885), .Z(net_11886) );
CLKBUF_X2 inst_17903 ( .A(net_17750), .Z(net_17751) );
CLKBUF_X2 inst_13728 ( .A(net_13575), .Z(net_13576) );
CLKBUF_X2 inst_13963 ( .A(net_13810), .Z(net_13811) );
CLKBUF_X2 inst_12410 ( .A(net_12257), .Z(net_12258) );
SDFF_X2 inst_1898 ( .D(net_7272), .SI(net_6969), .Q(net_6969), .SE(net_6283), .CK(net_14088) );
CLKBUF_X2 inst_15644 ( .A(net_14269), .Z(net_15492) );
INV_X2 inst_6275 ( .ZN(net_4326), .A(net_4276) );
SDFF_X2 inst_1714 ( .SI(net_7848), .Q(net_7848), .D(net_2702), .SE(net_2558), .CK(net_15250) );
AOI22_X2 inst_8551 ( .B2(net_4889), .A1(net_4803), .ZN(net_3240), .B1(net_3239), .A2(net_3097) );
AND2_X2 inst_9164 ( .A2(net_6105), .ZN(net_2864), .A1(net_2663) );
CLKBUF_X2 inst_14630 ( .A(net_14477), .Z(net_14478) );
CLKBUF_X2 inst_9428 ( .A(net_9258), .Z(net_9276) );
NAND2_X2 inst_4777 ( .ZN(net_1616), .A1(net_1615), .A2(net_1327) );
CLKBUF_X2 inst_15789 ( .A(net_15636), .Z(net_15637) );
CLKBUF_X2 inst_10762 ( .A(net_10609), .Z(net_10610) );
CLKBUF_X2 inst_10851 ( .A(net_10698), .Z(net_10699) );
CLKBUF_X2 inst_15333 ( .A(net_15180), .Z(net_15181) );
SDFF_X2 inst_1496 ( .SI(net_7853), .Q(net_7853), .D(net_2720), .SE(net_2558), .CK(net_18394) );
CLKBUF_X2 inst_11292 ( .A(net_11139), .Z(net_11140) );
AND2_X4 inst_9091 ( .ZN(net_2707), .A2(net_2381), .A1(net_2274) );
NAND2_X2 inst_4297 ( .A1(net_7091), .A2(net_5164), .ZN(net_5160) );
CLKBUF_X2 inst_9381 ( .A(net_9228), .Z(net_9229) );
CLKBUF_X2 inst_13005 ( .A(net_12136), .Z(net_12853) );
SDFF_X2 inst_1565 ( .Q(net_8041), .D(net_8041), .SI(net_2716), .SE(net_2545), .CK(net_17070) );
SDFF_X2 inst_924 ( .SI(net_8712), .Q(net_8712), .SE(net_6195), .D(net_3937), .CK(net_13015) );
XNOR2_X2 inst_287 ( .ZN(net_1008), .B(net_1007), .A(net_579) );
CLKBUF_X2 inst_10614 ( .A(net_10461), .Z(net_10462) );
AOI22_X2 inst_7929 ( .B1(net_8010), .A1(net_7976), .B2(net_6102), .A2(net_6097), .ZN(net_4195) );
CLKBUF_X2 inst_16144 ( .A(net_10999), .Z(net_15992) );
CLKBUF_X2 inst_12030 ( .A(net_11877), .Z(net_11878) );
OAI21_X2 inst_3094 ( .B1(net_2861), .ZN(net_2859), .B2(net_2491), .A(net_1836) );
CLKBUF_X2 inst_16305 ( .A(net_16152), .Z(net_16153) );
OAI33_X1 inst_2903 ( .ZN(net_3300), .B2(net_3299), .A3(net_3299), .A1(net_3246), .A2(net_2520), .B3(net_1306), .B1(net_1255) );
CLKBUF_X2 inst_13830 ( .A(net_10051), .Z(net_13678) );
NAND2_X4 inst_4045 ( .ZN(net_2559), .A1(net_2269), .A2(net_2267) );
CLKBUF_X2 inst_16749 ( .A(net_16596), .Z(net_16597) );
CLKBUF_X2 inst_12623 ( .A(net_12470), .Z(net_12471) );
NAND2_X2 inst_4890 ( .A2(net_7385), .ZN(net_706), .A1(net_174) );
SDFF_X2 inst_984 ( .D(net_7311), .SI(net_6619), .Q(net_6619), .SE(net_3123), .CK(net_9943) );
DFF_X1 inst_6734 ( .Q(net_6779), .D(net_5635), .CK(net_9206) );
SDFFS_X2 inst_2064 ( .SI(net_7396), .SE(net_2417), .Q(net_185), .D(net_185), .CK(net_14734), .SN(x6501) );
CLKBUF_X2 inst_14604 ( .A(net_11053), .Z(net_14452) );
CLKBUF_X2 inst_18546 ( .A(net_14292), .Z(net_18394) );
CLKBUF_X2 inst_15057 ( .A(net_12236), .Z(net_14905) );
SDFF_X2 inst_1292 ( .Q(net_8092), .D(net_8092), .SE(net_2707), .SI(net_2589), .CK(net_18411) );
CLKBUF_X2 inst_15769 ( .A(net_14541), .Z(net_15617) );
INV_X8 inst_5014 ( .ZN(net_4881), .A(net_4392) );
SDFF_X2 inst_1963 ( .D(net_7301), .SI(net_6958), .Q(net_6958), .SE(net_6281), .CK(net_15866) );
SDFF_X2 inst_1056 ( .SI(net_7321), .Q(net_6662), .D(net_6662), .SE(net_3126), .CK(net_9155) );
CLKBUF_X2 inst_11818 ( .A(net_11665), .Z(net_11666) );
CLKBUF_X2 inst_18611 ( .A(net_18458), .Z(net_18459) );
CLKBUF_X2 inst_17401 ( .A(net_17248), .Z(net_17249) );
NAND2_X2 inst_4247 ( .A1(net_6906), .A2(net_5247), .ZN(net_5213) );
NAND4_X2 inst_3648 ( .ZN(net_4913), .A3(net_4650), .A2(net_4519), .A4(net_4517), .A1(net_4458) );
CLKBUF_X2 inst_14434 ( .A(net_12143), .Z(net_14282) );
CLKBUF_X2 inst_14359 ( .A(net_11433), .Z(net_14207) );
INV_X2 inst_6524 ( .A(net_7431), .ZN(net_528) );
MUX2_X2 inst_4988 ( .A(net_9025), .Z(net_3960), .B(net_2818), .S(net_622) );
CLKBUF_X2 inst_11325 ( .A(net_11172), .Z(net_11173) );
CLKBUF_X2 inst_15074 ( .A(net_14921), .Z(net_14922) );
CLKBUF_X2 inst_14216 ( .A(net_12729), .Z(net_14064) );
CLKBUF_X2 inst_17815 ( .A(net_10292), .Z(net_17663) );
CLKBUF_X2 inst_11677 ( .A(net_10232), .Z(net_11525) );
CLKBUF_X2 inst_14996 ( .A(net_14843), .Z(net_14844) );
CLKBUF_X2 inst_18170 ( .A(net_16146), .Z(net_18018) );
CLKBUF_X2 inst_11559 ( .A(net_9580), .Z(net_11407) );
CLKBUF_X2 inst_10064 ( .A(net_9911), .Z(net_9912) );
CLKBUF_X2 inst_10999 ( .A(net_10846), .Z(net_10847) );
AND2_X4 inst_9077 ( .A1(net_6150), .ZN(net_3208), .A2(net_3072) );
AND4_X4 inst_9023 ( .ZN(net_5283), .A4(net_4865), .A3(net_4563), .A1(net_4556), .A2(net_4516) );
CLKBUF_X2 inst_10244 ( .A(net_10091), .Z(net_10092) );
CLKBUF_X2 inst_12714 ( .A(net_12094), .Z(net_12562) );
CLKBUF_X2 inst_14750 ( .A(net_14597), .Z(net_14598) );
CLKBUF_X2 inst_17876 ( .A(net_17723), .Z(net_17724) );
AOI22_X2 inst_8296 ( .B1(net_8694), .A1(net_8657), .B2(net_6109), .A2(net_3857), .ZN(net_3746) );
CLKBUF_X2 inst_12160 ( .A(net_12007), .Z(net_12008) );
CLKBUF_X2 inst_12246 ( .A(net_12093), .Z(net_12094) );
SDFF_X2 inst_1590 ( .Q(net_8019), .D(net_8019), .SI(net_2573), .SE(net_2545), .CK(net_15265) );
CLKBUF_X2 inst_17353 ( .A(net_12775), .Z(net_17201) );
INV_X2 inst_6229 ( .ZN(net_5481), .A(net_5310) );
CLKBUF_X2 inst_10648 ( .A(net_10495), .Z(net_10496) );
CLKBUF_X2 inst_10931 ( .A(net_10615), .Z(net_10779) );
CLKBUF_X2 inst_18093 ( .A(net_17940), .Z(net_17941) );
INV_X4 inst_5347 ( .ZN(net_2133), .A(net_1475) );
SDFFR_X2 inst_2318 ( .SE(net_2260), .Q(net_379), .D(net_379), .CK(net_11402), .RN(x6501), .SI(x1340) );
SDFF_X2 inst_399 ( .SI(net_8311), .Q(net_8311), .SE(net_3978), .D(net_3959), .CK(net_13212) );
CLKBUF_X2 inst_12433 ( .A(net_12280), .Z(net_12281) );
NAND3_X2 inst_3957 ( .A1(net_3046), .ZN(net_3039), .A3(net_3038), .A2(x2355) );
NAND2_X4 inst_4020 ( .A1(net_6147), .A2(net_6093), .ZN(net_4269) );
CLKBUF_X2 inst_9953 ( .A(net_9800), .Z(net_9801) );
CLKBUF_X2 inst_13404 ( .A(net_11836), .Z(net_13252) );
CLKBUF_X2 inst_17014 ( .A(net_16861), .Z(net_16862) );
SDFF_X2 inst_1299 ( .Q(net_8093), .D(net_8093), .SE(net_2707), .SI(net_2576), .CK(net_16085) );
INV_X2 inst_6450 ( .A(net_6326), .ZN(net_592) );
AOI22_X2 inst_8404 ( .B1(net_8749), .A1(net_8379), .A2(net_3867), .B2(net_3866), .ZN(net_3648) );
CLKBUF_X2 inst_10404 ( .A(net_10251), .Z(net_10252) );
CLKBUF_X2 inst_13487 ( .A(net_13334), .Z(net_13335) );
CLKBUF_X2 inst_17133 ( .A(net_16980), .Z(net_16981) );
SDFF_X2 inst_674 ( .Q(net_8413), .D(net_8413), .SI(net_3965), .SE(net_3934), .CK(net_10751) );
CLKBUF_X2 inst_14683 ( .A(net_14530), .Z(net_14531) );
INV_X4 inst_5259 ( .ZN(net_2073), .A(net_1885) );
INV_X4 inst_5518 ( .A(net_1575), .ZN(net_675) );
CLKBUF_X2 inst_14151 ( .A(net_13998), .Z(net_13999) );
CLKBUF_X2 inst_10859 ( .A(net_9116), .Z(net_10707) );
SDFFR_X2 inst_2253 ( .D(net_7394), .SE(net_2801), .SI(net_203), .Q(net_203), .CK(net_17772), .RN(x6501) );
CLKBUF_X2 inst_13670 ( .A(net_13517), .Z(net_13518) );
CLKBUF_X2 inst_18148 ( .A(net_17995), .Z(net_17996) );
CLKBUF_X2 inst_10115 ( .A(net_9962), .Z(net_9963) );
CLKBUF_X2 inst_9674 ( .A(net_9521), .Z(net_9522) );
CLKBUF_X2 inst_16255 ( .A(net_14249), .Z(net_16103) );
OR2_X2 inst_2868 ( .ZN(net_5727), .A2(net_5712), .A1(net_5679) );
INV_X2 inst_6522 ( .A(net_8900), .ZN(net_2101) );
CLKBUF_X2 inst_12254 ( .A(net_12101), .Z(net_12102) );
CLKBUF_X2 inst_18031 ( .A(net_14328), .Z(net_17879) );
CLKBUF_X2 inst_14549 ( .A(net_14396), .Z(net_14397) );
CLKBUF_X2 inst_12261 ( .A(net_9397), .Z(net_12109) );
SDFF_X2 inst_1832 ( .D(net_7298), .SI(net_6875), .Q(net_6875), .SE(net_6282), .CK(net_18188) );
CLKBUF_X2 inst_13241 ( .A(net_13088), .Z(net_13089) );
NAND2_X2 inst_4562 ( .ZN(net_3186), .A2(net_3185), .A1(net_3079) );
SDFF_X2 inst_640 ( .SI(net_8555), .Q(net_8555), .SE(net_3979), .D(net_3948), .CK(net_13477) );
CLKBUF_X2 inst_15740 ( .A(net_15587), .Z(net_15588) );
CLKBUF_X2 inst_9893 ( .A(net_9740), .Z(net_9741) );
DFFR_X1 inst_7500 ( .D(net_2388), .CK(net_13894), .RN(x6501), .Q(x661) );
CLKBUF_X2 inst_17785 ( .A(net_10561), .Z(net_17633) );
CLKBUF_X2 inst_16932 ( .A(net_16779), .Z(net_16780) );
SDFF_X2 inst_1478 ( .SI(net_7274), .Q(net_7091), .D(net_7091), .SE(net_6278), .CK(net_14133) );
INV_X4 inst_6098 ( .A(net_7258), .ZN(net_769) );
CLKBUF_X2 inst_18500 ( .A(net_17786), .Z(net_18348) );
CLKBUF_X2 inst_9535 ( .A(net_9382), .Z(net_9383) );
CLKBUF_X2 inst_17717 ( .A(net_17564), .Z(net_17565) );
AND2_X4 inst_9085 ( .A1(net_7628), .A2(net_2775), .ZN(net_2774) );
CLKBUF_X2 inst_12957 ( .A(net_12804), .Z(net_12805) );
CLKBUF_X2 inst_16661 ( .A(net_16035), .Z(net_16509) );
INV_X4 inst_6075 ( .A(net_7501), .ZN(net_3111) );
CLKBUF_X2 inst_13739 ( .A(net_10391), .Z(net_13587) );
CLKBUF_X2 inst_16977 ( .A(net_13018), .Z(net_16825) );
CLKBUF_X2 inst_16742 ( .A(net_16589), .Z(net_16590) );
SDFFS_X2 inst_2089 ( .SI(net_6831), .Q(net_6831), .D(net_6828), .SE(net_2146), .CK(net_18679), .SN(x6501) );
CLKBUF_X2 inst_15128 ( .A(net_14975), .Z(net_14976) );
CLKBUF_X2 inst_11378 ( .A(net_11225), .Z(net_11226) );
CLKBUF_X2 inst_16775 ( .A(net_16622), .Z(net_16623) );
SDFF_X2 inst_1679 ( .Q(net_8012), .D(net_8012), .SI(net_2705), .SE(net_2545), .CK(net_18529) );
CLKBUF_X2 inst_16280 ( .A(net_16127), .Z(net_16128) );
SDFFR_X2 inst_2215 ( .SI(net_2672), .SE(net_2477), .Q(net_305), .D(net_305), .CK(net_14719), .RN(x6501) );
SDFF_X2 inst_1855 ( .D(net_7264), .SI(net_6921), .Q(net_6921), .SE(net_6281), .CK(net_17418) );
XNOR2_X2 inst_337 ( .B(net_7389), .A(net_6371), .ZN(net_785) );
CLKBUF_X2 inst_11564 ( .A(net_11411), .Z(net_11412) );
CLKBUF_X2 inst_16575 ( .A(net_16212), .Z(net_16423) );
CLKBUF_X2 inst_11193 ( .A(net_11040), .Z(net_11041) );
INV_X2 inst_6220 ( .ZN(net_5490), .A(net_5349) );
CLKBUF_X2 inst_15355 ( .A(net_15202), .Z(net_15203) );
CLKBUF_X2 inst_13355 ( .A(net_13202), .Z(net_13203) );
CLKBUF_X2 inst_13775 ( .A(net_13622), .Z(net_13623) );
CLKBUF_X2 inst_9262 ( .A(net_9091), .Z(net_9110) );
CLKBUF_X2 inst_17249 ( .A(net_12326), .Z(net_17097) );
AOI22_X4 inst_7738 ( .A1(net_3292), .ZN(net_3176), .B1(net_3033), .B2(net_3032), .A2(net_2999) );
CLKBUF_X2 inst_18278 ( .A(net_18125), .Z(net_18126) );
SDFFR_X2 inst_2396 ( .SI(net_7374), .SE(net_2723), .D(net_2700), .QN(net_155), .CK(net_17812), .RN(x6501) );
CLKBUF_X2 inst_10232 ( .A(net_10079), .Z(net_10080) );
CLKBUF_X2 inst_15704 ( .A(net_15551), .Z(net_15552) );
CLKBUF_X2 inst_10281 ( .A(net_10128), .Z(net_10129) );
CLKBUF_X2 inst_14295 ( .A(net_14142), .Z(net_14143) );
CLKBUF_X2 inst_18589 ( .A(net_18436), .Z(net_18437) );
CLKBUF_X2 inst_14628 ( .A(net_14475), .Z(net_14476) );
INV_X4 inst_5908 ( .A(net_6301), .ZN(net_2688) );
XNOR2_X2 inst_246 ( .B(net_3029), .ZN(net_1212), .A(net_1211) );
NAND2_X2 inst_4443 ( .A1(net_6843), .A2(net_5016), .ZN(net_4984) );
SDFF_X2 inst_635 ( .SI(net_8549), .Q(net_8549), .SE(net_3979), .D(net_3940), .CK(net_10357) );
CLKBUF_X2 inst_12384 ( .A(net_12231), .Z(net_12232) );
INV_X4 inst_5787 ( .A(net_7637), .ZN(net_1459) );
AOI22_X2 inst_8510 ( .B1(net_6682), .A1(net_6649), .A2(net_6213), .B2(net_6138), .ZN(net_3430) );
CLKBUF_X2 inst_10569 ( .A(net_10416), .Z(net_10417) );
CLKBUF_X2 inst_16208 ( .A(net_16055), .Z(net_16056) );
CLKBUF_X2 inst_15140 ( .A(net_14987), .Z(net_14988) );
SDFF_X2 inst_519 ( .Q(net_8873), .D(net_8873), .SI(net_3956), .SE(net_3936), .CK(net_11018) );
NAND4_X2 inst_3796 ( .ZN(net_3630), .A1(net_3504), .A2(net_3503), .A3(net_3502), .A4(net_3501) );
CLKBUF_X2 inst_9359 ( .A(net_9156), .Z(net_9207) );
CLKBUF_X2 inst_12758 ( .A(net_12605), .Z(net_12606) );
CLKBUF_X2 inst_18198 ( .A(net_18045), .Z(net_18046) );
CLKBUF_X2 inst_12174 ( .A(net_12021), .Z(net_12022) );
SDFF_X2 inst_1053 ( .SI(net_7329), .Q(net_6670), .D(net_6670), .SE(net_3126), .CK(net_9515) );
INV_X4 inst_5158 ( .ZN(net_3295), .A(net_3122) );
DFFR_X2 inst_7231 ( .QN(net_6837), .D(net_2285), .CK(net_18728), .RN(x6501) );
CLKBUF_X2 inst_17639 ( .A(net_15404), .Z(net_17487) );
SDFFR_X1 inst_2774 ( .D(net_7387), .Q(net_7284), .SI(net_1957), .SE(net_1327), .CK(net_15378), .RN(x6501) );
CLKBUF_X2 inst_14673 ( .A(net_14520), .Z(net_14521) );
CLKBUF_X2 inst_17630 ( .A(net_17477), .Z(net_17478) );
DFFS_X2 inst_6871 ( .Q(net_8896), .D(net_4223), .CK(net_10680), .SN(x6501) );
CLKBUF_X2 inst_12202 ( .A(net_12049), .Z(net_12050) );
NAND2_X2 inst_4577 ( .ZN(net_6083), .A2(net_2996), .A1(net_2989) );
XNOR2_X2 inst_239 ( .ZN(net_1227), .A(net_1226), .B(net_1225) );
CLKBUF_X2 inst_18449 ( .A(net_18296), .Z(net_18297) );
CLKBUF_X2 inst_18098 ( .A(net_17945), .Z(net_17946) );
SDFF_X2 inst_1193 ( .D(net_7324), .SI(net_6566), .Q(net_6566), .SE(net_3070), .CK(net_12065) );
CLKBUF_X2 inst_14770 ( .A(net_14617), .Z(net_14618) );
CLKBUF_X2 inst_17703 ( .A(net_17550), .Z(net_17551) );
CLKBUF_X2 inst_18248 ( .A(net_18095), .Z(net_18096) );
CLKBUF_X2 inst_10582 ( .A(net_10429), .Z(net_10430) );
CLKBUF_X2 inst_15228 ( .A(net_15075), .Z(net_15076) );
CLKBUF_X2 inst_12395 ( .A(net_12242), .Z(net_12243) );
INV_X4 inst_6091 ( .A(net_6317), .ZN(net_1252) );
SDFF_X2 inst_601 ( .SI(net_8394), .Q(net_8394), .SE(net_3969), .D(net_3942), .CK(net_12613) );
DFFR_X1 inst_7391 ( .QN(net_6298), .D(net_5856), .CK(net_16780), .RN(x6501) );
CLKBUF_X2 inst_13709 ( .A(net_12008), .Z(net_13557) );
CLKBUF_X2 inst_18852 ( .A(net_18699), .Z(net_18700) );
AOI22_X2 inst_7952 ( .B1(net_8023), .A1(net_7989), .B2(net_6102), .A2(net_6097), .ZN(net_6034) );
AOI22_X2 inst_8097 ( .B1(net_8177), .A1(net_7735), .B2(net_6101), .A2(net_6095), .ZN(net_4050) );
SDFF_X2 inst_1773 ( .SI(net_8044), .Q(net_8044), .D(net_2721), .SE(net_2508), .CK(net_15733) );
CLKBUF_X2 inst_10133 ( .A(net_9948), .Z(net_9981) );
CLKBUF_X2 inst_10278 ( .A(net_10125), .Z(net_10126) );
SDFF_X2 inst_1583 ( .Q(net_8037), .D(net_8037), .SI(net_2639), .SE(net_2545), .CK(net_16489) );
SDFF_X2 inst_771 ( .Q(net_8781), .D(net_8781), .SI(net_3977), .SE(net_3879), .CK(net_11055) );
INV_X2 inst_6325 ( .ZN(net_3538), .A(net_3537) );
CLKBUF_X2 inst_11552 ( .A(net_9570), .Z(net_11400) );
CLKBUF_X2 inst_16002 ( .A(net_15849), .Z(net_15850) );
CLKBUF_X2 inst_15654 ( .A(net_11128), .Z(net_15502) );
DFFR_X2 inst_7324 ( .QN(net_395), .D(net_393), .CK(net_10805), .RN(x6501) );
DFFR_X1 inst_7402 ( .D(net_5743), .CK(net_16769), .RN(x6501), .Q(x468) );
CLKBUF_X2 inst_9334 ( .A(net_9159), .Z(net_9182) );
AOI22_X2 inst_8169 ( .A1(net_8603), .B1(net_8418), .ZN(net_3865), .A2(net_3864), .B2(net_3863) );
DFFR_X2 inst_7138 ( .QN(net_6402), .D(net_2928), .CK(net_17939), .RN(x6501) );
CLKBUF_X2 inst_12945 ( .A(net_10165), .Z(net_12793) );
INV_X4 inst_5782 ( .A(net_7599), .ZN(net_1093) );
CLKBUF_X2 inst_13873 ( .A(net_13720), .Z(net_13721) );
CLKBUF_X2 inst_10520 ( .A(net_10367), .Z(net_10368) );
SDFF_X2 inst_1319 ( .SI(net_7684), .Q(net_7684), .SE(net_2714), .D(net_2589), .CK(net_15627) );
SDFF_X2 inst_358 ( .Q(net_8756), .D(net_8756), .SE(net_3982), .SI(net_3973), .CK(net_10858) );
NAND2_X2 inst_4462 ( .ZN(net_4825), .A2(net_4660), .A1(net_4462) );
SDFF_X2 inst_1756 ( .Q(net_8209), .D(net_8209), .SI(net_2660), .SE(net_2561), .CK(net_16979) );
CLKBUF_X2 inst_14037 ( .A(net_13087), .Z(net_13885) );
CLKBUF_X2 inst_17041 ( .A(net_16888), .Z(net_16889) );
DFF_X1 inst_6766 ( .Q(net_7546), .D(net_4606), .CK(net_9720) );
AOI221_X2 inst_8794 ( .B2(net_5520), .C2(net_4965), .ZN(net_4903), .A(net_4641), .B1(net_283), .C1(net_274) );
DFFR_X2 inst_7108 ( .Q(net_8893), .D(net_3156), .CK(net_15695), .RN(x6501) );
CLKBUF_X2 inst_9309 ( .A(net_9156), .Z(net_9157) );
CLKBUF_X2 inst_15215 ( .A(net_15062), .Z(net_15063) );
CLKBUF_X2 inst_14177 ( .A(net_14024), .Z(net_14025) );
SDFF_X2 inst_655 ( .Q(net_8409), .D(net_8409), .SI(net_3943), .SE(net_3934), .CK(net_13108) );
INV_X4 inst_5914 ( .A(net_6373), .ZN(net_531) );
INV_X4 inst_5817 ( .A(net_6484), .ZN(net_1641) );
INV_X4 inst_5934 ( .A(net_6818), .ZN(net_4617) );
AOI22_X2 inst_8422 ( .B1(net_6662), .A1(net_6629), .A2(net_6213), .B2(net_6138), .ZN(net_3519) );
CLKBUF_X2 inst_9373 ( .A(net_9220), .Z(net_9221) );
CLKBUF_X2 inst_11316 ( .A(net_11163), .Z(net_11164) );
NAND2_X2 inst_4438 ( .A1(net_6875), .A2(net_5016), .ZN(net_4989) );
HA_X1 inst_6662 ( .S(net_3580), .CO(net_3579), .B(net_3265), .A(x2494) );
AOI221_X2 inst_8800 ( .B1(net_7184), .C2(net_6435), .B2(net_5655), .C1(net_5654), .ZN(net_4872), .A(net_4637) );
INV_X2 inst_6303 ( .ZN(net_3972), .A(net_3882) );
INV_X4 inst_5623 ( .A(net_7234), .ZN(net_1808) );
CLKBUF_X2 inst_9669 ( .A(net_9516), .Z(net_9517) );
CLKBUF_X2 inst_11996 ( .A(net_11843), .Z(net_11844) );
XOR2_X2 inst_41 ( .A(net_2921), .Z(net_1046), .B(net_514) );
CLKBUF_X2 inst_11516 ( .A(net_11363), .Z(net_11364) );
CLKBUF_X2 inst_11743 ( .A(net_11590), .Z(net_11591) );
CLKBUF_X2 inst_12569 ( .A(net_9410), .Z(net_12417) );
CLKBUF_X2 inst_18445 ( .A(net_18292), .Z(net_18293) );
SDFF_X2 inst_1989 ( .D(net_7277), .SI(net_7014), .Q(net_7014), .SE(net_6277), .CK(net_17332) );
CLKBUF_X2 inst_11868 ( .A(net_11715), .Z(net_11716) );
CLKBUF_X2 inst_13260 ( .A(net_13107), .Z(net_13108) );
XNOR2_X2 inst_152 ( .ZN(net_2036), .B(net_1930), .A(net_1929) );
CLKBUF_X2 inst_9694 ( .A(net_9431), .Z(net_9542) );
INV_X4 inst_5609 ( .A(net_8904), .ZN(net_1716) );
CLKBUF_X2 inst_11111 ( .A(net_10958), .Z(net_10959) );
DFFS_X1 inst_6944 ( .D(net_6145), .CK(net_13634), .SN(x6501), .Q(x757) );
CLKBUF_X2 inst_12314 ( .A(net_12042), .Z(net_12162) );
CLKBUF_X2 inst_18763 ( .A(net_12645), .Z(net_18611) );
INV_X2 inst_6388 ( .A(net_1352), .ZN(net_1300) );
SDFF_X2 inst_1400 ( .Q(net_8180), .D(net_8180), .SI(net_2721), .SE(net_2561), .CK(net_15848) );
CLKBUF_X2 inst_14374 ( .A(net_14221), .Z(net_14222) );
INV_X4 inst_5233 ( .ZN(net_2313), .A(net_2220) );
XOR2_X1 inst_89 ( .Z(net_1674), .B(net_1673), .A(net_1319) );
SDFF_X2 inst_1520 ( .Q(net_7889), .D(net_7889), .SI(net_2576), .SE(net_2543), .CK(net_16056) );
SDFF_X2 inst_1535 ( .Q(net_7986), .D(net_7986), .SI(net_2584), .SE(net_2542), .CK(net_15594) );
CLKBUF_X2 inst_13609 ( .A(net_13456), .Z(net_13457) );
CLKBUF_X2 inst_14112 ( .A(net_13959), .Z(net_13960) );
SDFF_X2 inst_788 ( .SI(net_8358), .Q(net_8358), .D(net_3955), .SE(net_3880), .CK(net_10516) );
CLKBUF_X2 inst_15525 ( .A(net_15372), .Z(net_15373) );
DFFR_X1 inst_7526 ( .D(net_6478), .Q(net_6475), .CK(net_11744), .RN(x6501) );
CLKBUF_X2 inst_13391 ( .A(net_12549), .Z(net_13239) );
CLKBUF_X2 inst_17174 ( .A(net_11646), .Z(net_17022) );
INV_X4 inst_5990 ( .A(net_7429), .ZN(net_3170) );
INV_X4 inst_5407 ( .A(net_8903), .ZN(net_1086) );
SDFF_X2 inst_1579 ( .Q(net_8030), .D(net_8030), .SI(net_2718), .SE(net_2545), .CK(net_15586) );
CLKBUF_X2 inst_13482 ( .A(net_13329), .Z(net_13330) );
XNOR2_X2 inst_193 ( .ZN(net_1552), .A(net_1116), .B(net_923) );
CLKBUF_X2 inst_14568 ( .A(net_9061), .Z(net_14416) );
CLKBUF_X2 inst_16153 ( .A(net_16000), .Z(net_16001) );
CLKBUF_X2 inst_17541 ( .A(net_17388), .Z(net_17389) );
CLKBUF_X2 inst_11704 ( .A(net_11551), .Z(net_11552) );
SDFF_X2 inst_1709 ( .Q(net_8018), .D(net_8018), .SI(net_2702), .SE(net_2545), .CK(net_15253) );
CLKBUF_X2 inst_16583 ( .A(net_16430), .Z(net_16431) );
CLKBUF_X2 inst_15358 ( .A(net_15205), .Z(net_15206) );
CLKBUF_X2 inst_17600 ( .A(net_17447), .Z(net_17448) );
DFFR_X1 inst_7531 ( .QN(net_6418), .D(net_1076), .CK(net_18015), .RN(x6501) );
SDFFR_X2 inst_2202 ( .QN(net_8905), .SE(net_6144), .D(net_2791), .SI(net_2790), .CK(net_17575), .RN(x6501) );
CLKBUF_X2 inst_11673 ( .A(net_11520), .Z(net_11521) );
OAI211_X2 inst_3180 ( .C2(net_6425), .ZN(net_5739), .A(net_5658), .C1(net_4950), .B(net_4827) );
AOI22_X2 inst_7969 ( .B1(net_7923), .A1(net_7821), .B2(net_6103), .A2(net_4398), .ZN(net_4160) );
NAND2_X2 inst_4737 ( .ZN(net_2711), .A2(net_1586), .A1(net_1361) );
CLKBUF_X2 inst_9965 ( .A(net_9812), .Z(net_9813) );
OAI21_X2 inst_2987 ( .B2(net_5912), .ZN(net_5909), .A(net_5802), .B1(net_733) );
CLKBUF_X2 inst_10618 ( .A(net_10465), .Z(net_10466) );
CLKBUF_X2 inst_15162 ( .A(net_15009), .Z(net_15010) );
CLKBUF_X2 inst_11645 ( .A(net_11492), .Z(net_11493) );
INV_X4 inst_5884 ( .A(net_7596), .ZN(net_1011) );
CLKBUF_X2 inst_11853 ( .A(net_11700), .Z(net_11701) );
CLKBUF_X2 inst_11170 ( .A(net_10742), .Z(net_11018) );
CLKBUF_X2 inst_12874 ( .A(net_12721), .Z(net_12722) );
SDFFR_X2 inst_2473 ( .D(net_7512), .SE(net_2313), .SI(net_428), .Q(net_428), .CK(net_14696), .RN(x6501) );
DFFR_X2 inst_7125 ( .QN(net_7354), .D(net_3062), .CK(net_9651), .RN(x6501) );
CLKBUF_X2 inst_17361 ( .A(net_10910), .Z(net_17209) );
NAND2_X2 inst_4516 ( .A2(net_6158), .ZN(net_3926), .A1(net_2887) );
CLKBUF_X2 inst_12442 ( .A(net_11513), .Z(net_12290) );
CLKBUF_X2 inst_13952 ( .A(net_10981), .Z(net_13800) );
OR2_X2 inst_2864 ( .ZN(net_5942), .A2(net_5941), .A1(net_2411) );
NOR2_X2 inst_3476 ( .ZN(net_2322), .A2(net_2166), .A1(net_1738) );
CLKBUF_X2 inst_14645 ( .A(net_14492), .Z(net_14493) );
NAND4_X2 inst_3789 ( .ZN(net_4232), .A1(net_3646), .A2(net_3645), .A3(net_3644), .A4(net_3643) );
CLKBUF_X2 inst_15001 ( .A(net_14848), .Z(net_14849) );
DFFR_X2 inst_7096 ( .QN(net_6471), .D(net_3343), .CK(net_15110), .RN(x6501) );
CLKBUF_X2 inst_16127 ( .A(net_12686), .Z(net_15975) );
SDFF_X2 inst_367 ( .SI(net_8552), .Q(net_8552), .SE(net_3979), .D(net_3976), .CK(net_12805) );
SDFF_X2 inst_957 ( .SI(net_7314), .Q(net_6688), .D(net_6688), .SE(net_3125), .CK(net_9950) );
CLKBUF_X2 inst_11589 ( .A(net_11436), .Z(net_11437) );
SDFF_X2 inst_1871 ( .D(net_7273), .SI(net_6970), .Q(net_6970), .SE(net_6283), .CK(net_14099) );
CLKBUF_X2 inst_16653 ( .A(net_16500), .Z(net_16501) );
INV_X2 inst_6460 ( .A(net_7217), .ZN(net_584) );
SDFFR_X2 inst_2300 ( .D(net_3205), .SE(net_2313), .SI(net_416), .Q(net_416), .CK(net_17293), .RN(x6501) );
DFFR_X1 inst_7552 ( .Q(net_7631), .D(net_1563), .CK(net_9816), .RN(x6501) );
CLKBUF_X2 inst_10800 ( .A(net_10647), .Z(net_10648) );
CLKBUF_X2 inst_18666 ( .A(net_18513), .Z(net_18514) );
SDFF_X2 inst_745 ( .Q(net_8801), .D(net_8801), .SI(net_3942), .SE(net_3879), .CK(net_10531) );
CLKBUF_X2 inst_11694 ( .A(net_11541), .Z(net_11542) );
DFFR_X2 inst_7024 ( .QN(net_6303), .D(net_5695), .CK(net_16932), .RN(x6501) );
CLKBUF_X2 inst_11622 ( .A(net_11469), .Z(net_11470) );
SDFF_X2 inst_2032 ( .SI(net_7776), .Q(net_7776), .D(net_2709), .SE(net_2459), .CK(net_15730) );
NAND2_X2 inst_4113 ( .ZN(net_5416), .A1(net_5143), .A2(net_5142) );
XOR2_X1 inst_80 ( .Z(net_3171), .B(net_3170), .A(net_3010) );
SDFF_X2 inst_836 ( .SI(net_8646), .Q(net_8646), .D(net_3944), .SE(net_3885), .CK(net_12250) );
AOI221_X2 inst_8821 ( .B1(net_8991), .C2(net_5538), .A(net_5520), .B2(net_5456), .ZN(net_4677), .C1(net_420) );
CLKBUF_X2 inst_9521 ( .A(net_9368), .Z(net_9369) );
INV_X2 inst_6564 ( .A(net_6373), .ZN(net_2148) );
CLKBUF_X2 inst_10771 ( .A(net_10618), .Z(net_10619) );
CLKBUF_X2 inst_9562 ( .A(net_9409), .Z(net_9410) );
XNOR2_X2 inst_241 ( .B(net_3330), .ZN(net_1220), .A(net_485) );
INV_X4 inst_5120 ( .ZN(net_4965), .A(net_4508) );
NAND2_X2 inst_4409 ( .A1(net_7049), .A2(net_5162), .ZN(net_5048) );
CLKBUF_X2 inst_16957 ( .A(net_16804), .Z(net_16805) );
MUX2_X2 inst_4934 ( .Z(net_3020), .A(net_3019), .B(net_3018), .S(x3712) );
CLKBUF_X2 inst_14705 ( .A(net_12290), .Z(net_14553) );
CLKBUF_X2 inst_16356 ( .A(net_11194), .Z(net_16204) );
CLKBUF_X2 inst_15384 ( .A(net_15231), .Z(net_15232) );
HA_X1 inst_6690 ( .S(net_2925), .CO(net_2924), .B(net_2915), .A(x2981) );
NAND3_X2 inst_3918 ( .ZN(net_5620), .A1(net_5549), .A3(net_5483), .A2(net_5319) );
CLKBUF_X2 inst_13491 ( .A(net_13338), .Z(net_13339) );
CLKBUF_X2 inst_14142 ( .A(net_11807), .Z(net_13990) );
CLKBUF_X2 inst_15534 ( .A(net_15381), .Z(net_15382) );
SDFFR_X1 inst_2758 ( .QN(net_7563), .D(net_3980), .SE(net_3144), .SI(net_2936), .CK(net_10879), .RN(x6501) );
NAND2_X2 inst_4504 ( .ZN(net_4367), .A2(net_4273), .A1(net_3926) );
SDFF_X2 inst_1116 ( .D(net_7320), .SI(net_6529), .Q(net_6529), .SE(net_3086), .CK(net_12078) );
AOI22_X2 inst_7947 ( .B1(net_8090), .A1(net_7750), .B2(net_6108), .A2(net_6096), .ZN(net_4179) );
CLKBUF_X2 inst_18311 ( .A(net_12984), .Z(net_18159) );
NAND4_X2 inst_3753 ( .ZN(net_4277), .A1(net_3996), .A2(net_3995), .A3(net_3994), .A4(net_3993) );
INV_X4 inst_5545 ( .ZN(net_879), .A(net_643) );
CLKBUF_X2 inst_12050 ( .A(net_11897), .Z(net_11898) );
CLKBUF_X2 inst_16393 ( .A(net_11934), .Z(net_16241) );
CLKBUF_X2 inst_17858 ( .A(net_11392), .Z(net_17706) );
CLKBUF_X2 inst_11555 ( .A(net_10517), .Z(net_11403) );
CLKBUF_X2 inst_17363 ( .A(net_17210), .Z(net_17211) );
INV_X2 inst_6394 ( .ZN(net_1174), .A(net_1173) );
OAI21_X2 inst_3136 ( .ZN(net_2064), .B2(net_2063), .A(net_2054), .B1(net_608) );
SDFF_X2 inst_402 ( .SI(net_8315), .Q(net_8315), .SE(net_3978), .D(net_3958), .CK(net_10036) );
CLKBUF_X2 inst_10962 ( .A(net_10809), .Z(net_10810) );
CLKBUF_X2 inst_16084 ( .A(net_15931), .Z(net_15932) );
CLKBUF_X2 inst_11259 ( .A(net_9686), .Z(net_11107) );
CLKBUF_X2 inst_13025 ( .A(net_12872), .Z(net_12873) );
INV_X4 inst_5832 ( .A(net_7437), .ZN(net_3390) );
CLKBUF_X2 inst_12815 ( .A(net_12662), .Z(net_12663) );
DFFR_X2 inst_7350 ( .Q(net_7340), .CK(net_11708), .D(x12915), .RN(x6501) );
SDFF_X2 inst_1288 ( .Q(net_7827), .D(net_7827), .SE(net_2730), .SI(net_2713), .CK(net_14441) );
NAND4_X2 inst_3844 ( .ZN(net_1720), .A1(net_1364), .A3(net_1027), .A2(net_1002), .A4(net_1001) );
CLKBUF_X2 inst_19128 ( .A(net_18975), .Z(net_18976) );
CLKBUF_X2 inst_11329 ( .A(net_11176), .Z(net_11177) );
SDFF_X2 inst_1033 ( .SI(net_7325), .Q(net_6732), .D(net_6732), .SE(net_3124), .CK(net_9139) );
CLKBUF_X2 inst_11845 ( .A(net_11344), .Z(net_11693) );
NAND2_X2 inst_4673 ( .ZN(net_2376), .A1(net_2115), .A2(net_2114) );
CLKBUF_X2 inst_14201 ( .A(net_14048), .Z(net_14049) );
CLKBUF_X2 inst_19081 ( .A(net_18928), .Z(net_18929) );
CLKBUF_X2 inst_16138 ( .A(net_15985), .Z(net_15986) );
INV_X4 inst_5582 ( .A(net_7357), .ZN(net_777) );
SDFF_X2 inst_1348 ( .Q(net_8203), .D(net_8203), .SI(net_2749), .SE(net_2561), .CK(net_14428) );
INV_X4 inst_5427 ( .ZN(net_2246), .A(net_834) );
SDFF_X2 inst_1748 ( .SI(net_7767), .Q(net_7767), .D(net_2660), .SE(net_2560), .CK(net_16984) );
CLKBUF_X2 inst_15686 ( .A(net_13684), .Z(net_15534) );
DFFR_X2 inst_7356 ( .Q(net_7334), .CK(net_11657), .D(x12969), .RN(x6501) );
CLKBUF_X2 inst_11423 ( .A(net_10998), .Z(net_11271) );
INV_X4 inst_5565 ( .ZN(net_1290), .A(net_665) );
CLKBUF_X2 inst_11684 ( .A(net_9571), .Z(net_11532) );
CLKBUF_X2 inst_14781 ( .A(net_14628), .Z(net_14629) );
CLKBUF_X2 inst_11864 ( .A(net_11711), .Z(net_11712) );
AOI222_X1 inst_8637 ( .C1(net_7442), .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_4213), .B1(net_3532), .A1(x13644) );
CLKBUF_X2 inst_9712 ( .A(net_9559), .Z(net_9560) );
CLKBUF_X2 inst_10145 ( .A(net_9992), .Z(net_9993) );
CLKBUF_X2 inst_14058 ( .A(net_13905), .Z(net_13906) );
CLKBUF_X2 inst_18211 ( .A(net_18058), .Z(net_18059) );
CLKBUF_X2 inst_9216 ( .A(net_9061), .Z(net_9064) );
CLKBUF_X2 inst_16439 ( .A(net_16286), .Z(net_16287) );
CLKBUF_X2 inst_19004 ( .A(net_18553), .Z(net_18852) );
CLKBUF_X2 inst_11088 ( .A(net_10935), .Z(net_10936) );
CLKBUF_X2 inst_12046 ( .A(net_10016), .Z(net_11894) );
INV_X2 inst_6397 ( .ZN(net_1163), .A(net_1162) );
DFFR_X2 inst_7337 ( .Q(net_7313), .CK(net_11390), .D(x13163), .RN(x6501) );
SDFFR_X2 inst_2461 ( .D(net_6321), .SE(net_2313), .SI(net_443), .Q(net_443), .CK(net_14698), .RN(x6501) );
CLKBUF_X2 inst_18420 ( .A(net_18267), .Z(net_18268) );
AOI221_X2 inst_8814 ( .C2(net_5535), .B2(net_5260), .A(net_4898), .ZN(net_4713), .B1(net_3544), .C1(net_457) );
SDFF_X2 inst_732 ( .SI(net_8370), .Q(net_8370), .D(net_3948), .SE(net_3880), .CK(net_13399) );
CLKBUF_X2 inst_12183 ( .A(net_12030), .Z(net_12031) );
CLKBUF_X2 inst_13044 ( .A(net_12891), .Z(net_12892) );
AOI22_X2 inst_8023 ( .B1(net_8066), .A1(net_7862), .B2(net_6107), .ZN(net_6016), .A2(net_4400) );
INV_X4 inst_5968 ( .A(net_7426), .ZN(net_2921) );
XOR2_X1 inst_79 ( .B(net_3334), .Z(net_3172), .A(net_3012) );
CLKBUF_X2 inst_11250 ( .A(net_11097), .Z(net_11098) );
AOI21_X2 inst_8930 ( .B2(net_5843), .ZN(net_5681), .A(net_5666), .B1(x364) );
SDFFR_X1 inst_2654 ( .D(net_6776), .SE(net_4506), .CK(net_9188), .RN(x6501), .SI(x1597), .Q(x1597) );
DFFR_X2 inst_7088 ( .QN(net_7347), .D(net_6158), .CK(net_9574), .RN(x6501) );
CLKBUF_X2 inst_16526 ( .A(net_12153), .Z(net_16374) );
CLKBUF_X2 inst_16691 ( .A(net_16538), .Z(net_16539) );
CLKBUF_X2 inst_11662 ( .A(net_11341), .Z(net_11510) );
AOI221_X2 inst_8838 ( .C1(net_8179), .B1(net_7737), .C2(net_6101), .B2(net_6095), .ZN(net_5993), .A(net_4284) );
CLKBUF_X2 inst_11962 ( .A(net_9659), .Z(net_11810) );
AOI22_X2 inst_7895 ( .B1(net_8977), .A2(net_5538), .B2(net_5456), .ZN(net_4534), .A1(net_406) );
NAND2_X2 inst_4413 ( .A1(net_6852), .A2(net_5016), .ZN(net_5014) );
CLKBUF_X2 inst_16293 ( .A(net_16140), .Z(net_16141) );
CLKBUF_X2 inst_17938 ( .A(net_17785), .Z(net_17786) );
OAI221_X2 inst_2975 ( .ZN(net_2208), .B1(net_2207), .C1(net_2206), .A(net_2011), .C2(net_2010), .B2(net_1925) );
SDFF_X2 inst_1741 ( .SI(net_7302), .Q(net_7079), .D(net_7079), .SE(net_6280), .CK(net_15432) );
INV_X4 inst_5594 ( .A(net_5967), .ZN(x3156) );
SDFF_X2 inst_1658 ( .SI(net_7748), .Q(net_7748), .D(net_2584), .SE(net_2560), .CK(net_18851) );
INV_X2 inst_6515 ( .ZN(net_905), .A(net_229) );
CLKBUF_X2 inst_14991 ( .A(net_14838), .Z(net_14839) );
AOI211_X2 inst_9003 ( .ZN(net_5713), .A(net_5590), .C2(net_5463), .B(net_4819), .C1(net_443) );
NAND2_X2 inst_4267 ( .A1(net_6915), .A2(net_5247), .ZN(net_5193) );
NAND3_X2 inst_3965 ( .A2(net_7645), .A1(net_6264), .A3(net_5691), .ZN(net_2452) );
CLKBUF_X2 inst_12829 ( .A(net_10386), .Z(net_12677) );
SDFF_X2 inst_440 ( .Q(net_8769), .D(net_8769), .SE(net_3982), .SI(net_3953), .CK(net_10293) );
CLKBUF_X2 inst_18963 ( .A(net_18810), .Z(net_18811) );
CLKBUF_X2 inst_14386 ( .A(net_11471), .Z(net_14234) );
MUX2_X2 inst_4927 ( .S(net_3552), .Z(net_3551), .A(net_3550), .B(net_1021) );
SDFF_X2 inst_1887 ( .D(net_7301), .SI(net_6998), .Q(net_6998), .SE(net_6283), .CK(net_15874) );
CLKBUF_X2 inst_15287 ( .A(net_15134), .Z(net_15135) );
CLKBUF_X2 inst_15423 ( .A(net_15270), .Z(net_15271) );
CLKBUF_X2 inst_11708 ( .A(net_11555), .Z(net_11556) );
CLKBUF_X2 inst_15108 ( .A(net_9959), .Z(net_14956) );
NOR2_X2 inst_3579 ( .ZN(net_1302), .A1(net_1092), .A2(net_1091) );
CLKBUF_X2 inst_16560 ( .A(net_16385), .Z(net_16408) );
CLKBUF_X2 inst_16537 ( .A(net_16384), .Z(net_16385) );
INV_X4 inst_5688 ( .ZN(net_1052), .A(net_148) );
SDFF_X2 inst_1672 ( .SI(net_7771), .Q(net_7771), .D(net_2703), .SE(net_2560), .CK(net_14001) );
CLKBUF_X2 inst_16921 ( .A(net_16768), .Z(net_16769) );
CLKBUF_X2 inst_13705 ( .A(net_12774), .Z(net_13553) );
AOI222_X1 inst_8625 ( .A2(net_8253), .B1(net_7595), .C2(net_6117), .ZN(net_4801), .A1(net_4800), .B2(net_4799), .C1(net_2666) );
CLKBUF_X2 inst_12120 ( .A(net_11967), .Z(net_11968) );
CLKBUF_X2 inst_17661 ( .A(net_12541), .Z(net_17509) );
SDFF_X2 inst_2015 ( .SI(net_7936), .Q(net_7936), .D(net_2715), .SE(net_2461), .CK(net_14153) );
CLKBUF_X2 inst_18110 ( .A(net_17957), .Z(net_17958) );
CLKBUF_X2 inst_12108 ( .A(net_11955), .Z(net_11956) );
NAND3_X2 inst_3937 ( .ZN(net_4940), .A1(net_4794), .A3(net_4710), .A2(net_4492) );
OAI221_X2 inst_2970 ( .B2(net_2489), .ZN(net_2455), .C2(net_2450), .A(net_2270), .B1(net_1934), .C1(net_674) );
CLKBUF_X2 inst_14488 ( .A(net_14335), .Z(net_14336) );
CLKBUF_X2 inst_11950 ( .A(net_10995), .Z(net_11798) );
CLKBUF_X2 inst_10942 ( .A(net_10789), .Z(net_10790) );
AOI22_X2 inst_8278 ( .B1(net_8766), .A1(net_8396), .A2(net_3867), .B2(net_3866), .ZN(net_3763) );
CLKBUF_X2 inst_9281 ( .A(net_9078), .Z(net_9129) );
NAND2_X2 inst_4085 ( .ZN(net_5756), .A1(net_5718), .A2(net_5599) );
CLKBUF_X2 inst_16360 ( .A(net_16207), .Z(net_16208) );
CLKBUF_X2 inst_18576 ( .A(net_18423), .Z(net_18424) );
CLKBUF_X2 inst_14719 ( .A(net_14566), .Z(net_14567) );
CLKBUF_X2 inst_18194 ( .A(net_18041), .Z(net_18042) );
CLKBUF_X2 inst_17058 ( .A(net_16905), .Z(net_16906) );
CLKBUF_X2 inst_13183 ( .A(net_9542), .Z(net_13031) );
MUX2_X2 inst_4990 ( .S(net_8901), .A(net_8250), .Z(net_2791), .B(net_1162) );
INV_X4 inst_5664 ( .ZN(net_1057), .A(x12810) );
CLKBUF_X2 inst_10317 ( .A(net_10164), .Z(net_10165) );
CLKBUF_X2 inst_12285 ( .A(net_10024), .Z(net_12133) );
CLKBUF_X2 inst_9442 ( .A(net_9289), .Z(net_9290) );
CLKBUF_X2 inst_11090 ( .A(net_10937), .Z(net_10938) );
SDFF_X2 inst_815 ( .SI(net_8506), .Q(net_8506), .D(net_3955), .SE(net_3884), .CK(net_13236) );
SDFFR_X2 inst_2165 ( .QN(net_7587), .D(net_3975), .SE(net_3144), .SI(net_3136), .CK(net_12652), .RN(x6501) );
CLKBUF_X2 inst_15433 ( .A(net_15280), .Z(net_15281) );
OAI21_X2 inst_3081 ( .A(net_3246), .ZN(net_3244), .B1(net_646), .B2(x13291) );
INV_X4 inst_5187 ( .A(net_4928), .ZN(net_4891) );
CLKBUF_X2 inst_12096 ( .A(net_10383), .Z(net_11944) );
AOI22_X2 inst_8227 ( .B1(net_8759), .A1(net_8389), .A2(net_3867), .B2(net_3866), .ZN(net_3810) );
CLKBUF_X2 inst_16330 ( .A(net_16177), .Z(net_16178) );
DFFR_X2 inst_7006 ( .QN(net_5973), .D(net_5840), .CK(net_11544), .RN(x6501) );
AOI21_X2 inst_8888 ( .B2(net_5871), .ZN(net_5810), .A(net_5809), .B1(net_2690) );
SDFFR_X2 inst_2108 ( .SI(net_7408), .Q(net_7408), .SE(net_6198), .D(net_5732), .CK(net_9380), .RN(x6501) );
NOR2_X2 inst_3572 ( .A1(net_7399), .ZN(net_4322), .A2(net_664) );
AOI22_X2 inst_7761 ( .B1(net_6989), .A1(net_6949), .A2(net_5443), .B2(net_5442), .ZN(net_5362) );
CLKBUF_X2 inst_12178 ( .A(net_12025), .Z(net_12026) );
CLKBUF_X2 inst_11177 ( .A(net_11024), .Z(net_11025) );
SDFF_X2 inst_413 ( .SI(net_8299), .Q(net_8299), .D(net_3980), .SE(net_3978), .CK(net_13366) );
INV_X4 inst_5094 ( .ZN(net_5703), .A(net_5678) );
AOI22_X2 inst_8118 ( .A1(net_7945), .B1(net_7775), .A2(net_6092), .B2(net_6091), .ZN(net_4030) );
INV_X16 inst_6623 ( .ZN(net_4816), .A(net_4708) );
SDFF_X2 inst_859 ( .Q(net_8566), .D(net_8566), .SI(net_3960), .SE(net_3878), .CK(net_13316) );
CLKBUF_X2 inst_13446 ( .A(net_13293), .Z(net_13294) );
NOR2_X4 inst_3323 ( .ZN(net_4962), .A1(net_4783), .A2(net_4557) );
CLKBUF_X2 inst_12634 ( .A(net_12481), .Z(net_12482) );
CLKBUF_X2 inst_17448 ( .A(net_17295), .Z(net_17296) );
CLKBUF_X2 inst_13013 ( .A(net_11201), .Z(net_12861) );
CLKBUF_X2 inst_18391 ( .A(net_18238), .Z(net_18239) );
INV_X4 inst_5938 ( .A(net_7255), .ZN(net_1953) );
CLKBUF_X2 inst_13061 ( .A(net_11653), .Z(net_12909) );
INV_X4 inst_5736 ( .A(net_8927), .ZN(net_4522) );
SDFF_X2 inst_1691 ( .SI(net_7861), .Q(net_7861), .D(net_2713), .SE(net_2558), .CK(net_13752) );
CLKBUF_X2 inst_15626 ( .A(net_15473), .Z(net_15474) );
AOI211_X2 inst_9019 ( .ZN(net_1919), .B(net_1658), .C2(net_1657), .A(net_1326), .C1(net_1325) );
CLKBUF_X2 inst_11156 ( .A(net_11003), .Z(net_11004) );
CLKBUF_X2 inst_15413 ( .A(net_9146), .Z(net_15261) );
NAND4_X2 inst_3688 ( .A4(net_6246), .A1(net_6245), .ZN(net_4449), .A2(net_3840), .A3(net_3839) );
INV_X4 inst_5476 ( .ZN(net_868), .A(net_744) );
INV_X4 inst_5776 ( .A(net_7507), .ZN(net_3203) );
CLKBUF_X2 inst_18863 ( .A(net_18710), .Z(net_18711) );
CLKBUF_X2 inst_12149 ( .A(net_9523), .Z(net_11997) );
CLKBUF_X2 inst_10186 ( .A(net_9932), .Z(net_10034) );
CLKBUF_X2 inst_13124 ( .A(net_12971), .Z(net_12972) );
SDFF_X2 inst_560 ( .Q(net_8675), .D(net_8675), .SI(net_3937), .SE(net_3935), .CK(net_12449) );
CLKBUF_X2 inst_11167 ( .A(net_11014), .Z(net_11015) );
INV_X4 inst_5393 ( .ZN(net_1081), .A(net_1080) );
INV_X4 inst_5199 ( .ZN(net_2586), .A(net_2470) );
CLKBUF_X2 inst_9729 ( .A(net_9576), .Z(net_9577) );
CLKBUF_X2 inst_12953 ( .A(net_12800), .Z(net_12801) );
DFFR_X1 inst_7479 ( .QN(net_7438), .D(net_4218), .CK(net_12851), .RN(x6501) );
NAND2_X2 inst_4809 ( .A1(net_9009), .A2(net_2429), .ZN(net_2233) );
SDFF_X2 inst_1802 ( .SI(net_8061), .Q(net_8061), .D(net_2719), .SE(net_2508), .CK(net_18755) );
CLKBUF_X2 inst_10260 ( .A(net_10107), .Z(net_10108) );
DFF_X1 inst_6851 ( .Q(net_6439), .D(net_3630), .CK(net_17896) );
OAI21_X4 inst_2982 ( .ZN(net_3180), .A(net_2995), .B2(net_2941), .B1(net_1211) );
CLKBUF_X2 inst_15444 ( .A(net_15291), .Z(net_15292) );
CLKBUF_X2 inst_11837 ( .A(net_11684), .Z(net_11685) );
NOR2_X2 inst_3359 ( .ZN(net_5566), .A1(net_5392), .A2(net_5391) );
CLKBUF_X2 inst_10100 ( .A(net_9078), .Z(net_9948) );
CLKBUF_X2 inst_18974 ( .A(net_13351), .Z(net_18822) );
DFFR_X1 inst_7491 ( .QN(net_6474), .D(net_3340), .CK(net_15141), .RN(x6501) );
CLKBUF_X2 inst_14338 ( .A(net_14185), .Z(net_14186) );
NAND2_X2 inst_4418 ( .A1(net_6857), .A2(net_5016), .ZN(net_5009) );
XOR2_X1 inst_96 ( .Z(net_1392), .B(net_1391), .A(net_705) );
NAND2_X2 inst_4346 ( .A1(net_7066), .A2(net_5162), .ZN(net_5111) );
AOI22_X2 inst_8564 ( .B1(net_2473), .ZN(net_2329), .A2(net_2328), .B2(net_2327), .A1(net_2248) );
CLKBUF_X2 inst_18705 ( .A(net_14156), .Z(net_18553) );
CLKBUF_X2 inst_17156 ( .A(net_17003), .Z(net_17004) );
CLKBUF_X2 inst_11205 ( .A(net_11052), .Z(net_11053) );
CLKBUF_X2 inst_9330 ( .A(net_9177), .Z(net_9178) );
CLKBUF_X2 inst_18687 ( .A(net_15224), .Z(net_18535) );
CLKBUF_X2 inst_17616 ( .A(net_17368), .Z(net_17464) );
CLKBUF_X2 inst_10912 ( .A(net_9983), .Z(net_10760) );
CLKBUF_X2 inst_15558 ( .A(net_15405), .Z(net_15406) );
CLKBUF_X2 inst_14575 ( .A(net_14422), .Z(net_14423) );
CLKBUF_X2 inst_15937 ( .A(net_15784), .Z(net_15785) );
SDFFR_X2 inst_2436 ( .D(net_3546), .SE(net_2313), .SI(net_430), .Q(net_430), .CK(net_16414), .RN(x6501) );
OR2_X4 inst_2832 ( .ZN(net_3144), .A2(net_2952), .A1(net_2233) );
CLKBUF_X2 inst_19168 ( .A(net_17819), .Z(net_19016) );
SDFF_X2 inst_603 ( .SI(net_8397), .Q(net_8397), .D(net_3975), .SE(net_3969), .CK(net_12540) );
XNOR2_X2 inst_291 ( .B(net_7382), .ZN(net_1001), .A(net_545) );
CLKBUF_X2 inst_9488 ( .A(net_9335), .Z(net_9336) );
CLKBUF_X2 inst_15521 ( .A(net_15368), .Z(net_15369) );
CLKBUF_X2 inst_12213 ( .A(net_9899), .Z(net_12061) );
CLKBUF_X2 inst_16569 ( .A(net_16416), .Z(net_16417) );
CLKBUF_X2 inst_18709 ( .A(net_18556), .Z(net_18557) );
CLKBUF_X2 inst_16846 ( .A(net_16693), .Z(net_16694) );
CLKBUF_X2 inst_16688 ( .A(net_16335), .Z(net_16536) );
DFF_X1 inst_6849 ( .Q(net_6437), .D(net_3632), .CK(net_17903) );
CLKBUF_X2 inst_10310 ( .A(net_9251), .Z(net_10158) );
AND2_X4 inst_9110 ( .ZN(net_2069), .A2(net_2046), .A1(net_1870) );
INV_X2 inst_6512 ( .A(net_6351), .ZN(net_2130) );
DFFS_X1 inst_6925 ( .D(net_6145), .CK(net_16373), .SN(x6501), .Q(x820) );
AOI22_X2 inst_7745 ( .B1(net_6974), .A1(net_6934), .A2(net_5443), .B2(net_5442), .ZN(net_5426) );
SDFF_X2 inst_1807 ( .SI(net_6956), .Q(net_6956), .SE(net_6281), .D(net_2544), .CK(net_15881) );
AOI222_X1 inst_8600 ( .A2(net_6757), .B2(net_6198), .A1(net_5835), .ZN(net_5825), .C2(net_5824), .C1(net_2079), .B1(net_1931) );
DFFR_X2 inst_7236 ( .QN(net_8217), .D(net_2178), .CK(net_17302), .RN(x6501) );
CLKBUF_X2 inst_9989 ( .A(net_9836), .Z(net_9837) );
SDFF_X2 inst_913 ( .SI(net_8733), .Q(net_8733), .SE(net_6195), .D(net_3952), .CK(net_10314) );
CLKBUF_X2 inst_12274 ( .A(net_12121), .Z(net_12122) );
CLKBUF_X2 inst_12712 ( .A(net_10289), .Z(net_12560) );
CLKBUF_X2 inst_18267 ( .A(net_14025), .Z(net_18115) );
CLKBUF_X2 inst_15999 ( .A(net_15846), .Z(net_15847) );
CLKBUF_X2 inst_16434 ( .A(net_16281), .Z(net_16282) );
CLKBUF_X2 inst_17567 ( .A(net_17414), .Z(net_17415) );
CLKBUF_X2 inst_18120 ( .A(net_9927), .Z(net_17968) );
CLKBUF_X2 inst_15188 ( .A(net_13860), .Z(net_15036) );
CLKBUF_X2 inst_15502 ( .A(net_15349), .Z(net_15350) );
INV_X16 inst_6633 ( .ZN(net_3866), .A(net_3366) );
CLKBUF_X2 inst_10322 ( .A(net_10169), .Z(net_10170) );
CLKBUF_X2 inst_12004 ( .A(net_11851), .Z(net_11852) );
CLKBUF_X2 inst_9298 ( .A(net_9145), .Z(net_9146) );
CLKBUF_X2 inst_11214 ( .A(net_11061), .Z(net_11062) );
SDFFR_X2 inst_2483 ( .Q(net_8982), .D(net_8982), .SI(net_4526), .SE(net_2562), .CK(net_16639), .RN(x6501) );
SDFF_X2 inst_1414 ( .SI(net_7286), .Q(net_7143), .D(net_7143), .SE(net_6279), .CK(net_16235) );
CLKBUF_X2 inst_16101 ( .A(net_15948), .Z(net_15949) );
CLKBUF_X2 inst_17658 ( .A(net_17505), .Z(net_17506) );
AOI22_X2 inst_8451 ( .B1(net_6603), .A1(net_6570), .A2(net_6257), .B2(net_6110), .ZN(net_3489) );
NAND3_X2 inst_3994 ( .A2(net_9006), .ZN(net_1928), .A1(net_1661), .A3(net_1179) );
SDFF_X2 inst_449 ( .Q(net_8746), .D(net_8746), .SE(net_3982), .SI(net_3965), .CK(net_10770) );
CLKBUF_X2 inst_10797 ( .A(net_10644), .Z(net_10645) );
CLKBUF_X2 inst_10354 ( .A(net_10201), .Z(net_10202) );
SDFFR_X1 inst_2790 ( .Q(net_7288), .D(net_2796), .SI(net_1954), .SE(net_1327), .CK(net_15361), .RN(x6501) );
SDFFR_X2 inst_2138 ( .SI(net_7178), .Q(net_7178), .D(net_6429), .SE(net_4362), .CK(net_13556), .RN(x6501) );
DFFR_X2 inst_7152 ( .QN(net_7517), .D(net_2826), .CK(net_17632), .RN(x6501) );
INV_X4 inst_5599 ( .A(net_7427), .ZN(net_3048) );
CLKBUF_X2 inst_16823 ( .A(net_16670), .Z(net_16671) );
INV_X2 inst_6593 ( .A(net_6126), .ZN(net_6125) );
CLKBUF_X2 inst_11417 ( .A(net_11264), .Z(net_11265) );
INV_X4 inst_6055 ( .A(net_6795), .ZN(net_1209) );
CLKBUF_X2 inst_13362 ( .A(net_13209), .Z(net_13210) );
NOR4_X2 inst_3249 ( .A1(net_2697), .A2(net_2696), .A3(net_2695), .ZN(net_1256), .A4(net_1052) );
MUX2_X2 inst_4935 ( .Z(net_2962), .S(net_2782), .A(net_2781), .B(net_2185) );
CLKBUF_X2 inst_17505 ( .A(net_12825), .Z(net_17353) );
AOI21_X2 inst_8961 ( .ZN(net_3586), .B2(net_3578), .B1(net_3035), .A(net_3027) );
DFFR_X1 inst_7498 ( .Q(net_6407), .D(net_2446), .CK(net_9678), .RN(x6501) );
CLKBUF_X2 inst_9860 ( .A(net_9299), .Z(net_9708) );
CLKBUF_X2 inst_12420 ( .A(net_12267), .Z(net_12268) );
CLKBUF_X2 inst_13369 ( .A(net_10441), .Z(net_13217) );
CLKBUF_X2 inst_11044 ( .A(net_10891), .Z(net_10892) );
CLKBUF_X2 inst_12973 ( .A(net_9114), .Z(net_12821) );
CLKBUF_X2 inst_19103 ( .A(net_18950), .Z(net_18951) );
AOI22_X2 inst_8201 ( .A1(net_8607), .B1(net_8422), .A2(net_3864), .B2(net_3863), .ZN(net_3835) );
NOR2_X2 inst_3614 ( .A2(net_7488), .A1(net_7487), .ZN(net_1099) );
AOI21_X2 inst_8893 ( .B2(net_5871), .ZN(net_5794), .A(net_5788), .B1(x451) );
CLKBUF_X2 inst_18672 ( .A(net_17144), .Z(net_18520) );
CLKBUF_X2 inst_16224 ( .A(net_16071), .Z(net_16072) );
CLKBUF_X2 inst_12776 ( .A(net_9991), .Z(net_12624) );
SDFF_X2 inst_588 ( .Q(net_8824), .D(net_8824), .SE(net_3964), .SI(net_3946), .CK(net_10727) );
CLKBUF_X2 inst_10752 ( .A(net_9300), .Z(net_10600) );
CLKBUF_X2 inst_10394 ( .A(net_10241), .Z(net_10242) );
CLKBUF_X2 inst_11411 ( .A(net_11258), .Z(net_11259) );
CLKBUF_X2 inst_16488 ( .A(net_16335), .Z(net_16336) );
CLKBUF_X2 inst_17296 ( .A(net_17143), .Z(net_17144) );
CLKBUF_X2 inst_14015 ( .A(net_13862), .Z(net_13863) );
CLKBUF_X2 inst_10329 ( .A(net_10176), .Z(net_10177) );
CLKBUF_X2 inst_9405 ( .A(net_9063), .Z(net_9253) );
CLKBUF_X2 inst_16557 ( .A(net_16404), .Z(net_16405) );
CLKBUF_X2 inst_19063 ( .A(net_18910), .Z(net_18911) );
CLKBUF_X2 inst_11060 ( .A(net_10907), .Z(net_10908) );
NAND2_X2 inst_4752 ( .ZN(net_2576), .A2(net_1586), .A1(net_1363) );
SDFF_X2 inst_1356 ( .Q(net_8190), .D(net_8190), .SI(net_2584), .SE(net_2561), .CK(net_15608) );
CLKBUF_X2 inst_12913 ( .A(net_12760), .Z(net_12761) );
INV_X2 inst_6447 ( .ZN(net_599), .A(x6501) );
SDFFR_X2 inst_2628 ( .Q(net_7388), .D(net_7388), .SE(net_1136), .CK(net_15864), .RN(x6501), .SI(x4570) );
SDFFR_X2 inst_2196 ( .D(net_2768), .SE(net_2519), .SI(net_303), .Q(net_303), .CK(net_13722), .RN(x6501) );
CLKBUF_X2 inst_14159 ( .A(net_13004), .Z(net_14007) );
AOI22_X2 inst_7754 ( .B1(net_6982), .A1(net_6942), .A2(net_5443), .B2(net_5442), .ZN(net_5390) );
DFFR_X2 inst_7145 ( .QN(net_6397), .D(net_2877), .CK(net_15685), .RN(x6501) );
CLKBUF_X2 inst_14083 ( .A(net_10521), .Z(net_13931) );
SDFF_X2 inst_1045 ( .SI(net_7328), .Q(net_6702), .D(net_6702), .SE(net_3125), .CK(net_9135) );
CLKBUF_X2 inst_18054 ( .A(net_17901), .Z(net_17902) );
CLKBUF_X2 inst_18042 ( .A(net_12853), .Z(net_17890) );
XNOR2_X2 inst_252 ( .A(net_6296), .B(net_2736), .ZN(net_1197) );
SDFF_X2 inst_865 ( .Q(net_8574), .D(net_8574), .SI(net_3958), .SE(net_3878), .CK(net_13159) );
SDFF_X2 inst_956 ( .SI(net_7310), .Q(net_6717), .D(net_6717), .SE(net_3125), .CK(net_11918) );
CLKBUF_X2 inst_10959 ( .A(net_10806), .Z(net_10807) );
CLKBUF_X2 inst_17269 ( .A(net_12699), .Z(net_17117) );
CLKBUF_X2 inst_18827 ( .A(net_18674), .Z(net_18675) );
CLKBUF_X2 inst_10177 ( .A(net_10024), .Z(net_10025) );
NAND2_X2 inst_4684 ( .A2(net_2282), .ZN(net_2199), .A1(net_2031) );
CLKBUF_X2 inst_12757 ( .A(net_12604), .Z(net_12605) );
SDFF_X2 inst_484 ( .SI(net_8607), .Q(net_8607), .SE(net_3984), .D(net_3959), .CK(net_10177) );
CLKBUF_X2 inst_16041 ( .A(net_10898), .Z(net_15889) );
NAND2_X2 inst_4474 ( .A2(net_5657), .ZN(net_4643), .A1(net_573) );
CLKBUF_X2 inst_9272 ( .A(net_9119), .Z(net_9120) );
CLKBUF_X2 inst_15902 ( .A(net_12001), .Z(net_15750) );
XOR2_X2 inst_32 ( .A(net_6485), .Z(net_1205), .B(net_589) );
AND2_X4 inst_9129 ( .ZN(net_1405), .A2(net_888), .A1(net_163) );
SDFF_X2 inst_1821 ( .D(net_7295), .SI(net_7032), .Q(net_7032), .SE(net_6277), .CK(net_15418) );
CLKBUF_X2 inst_16316 ( .A(net_16163), .Z(net_16164) );
DFFR_X2 inst_7271 ( .Q(net_5955), .D(net_2009), .CK(net_11811), .RN(x6501) );
SDFF_X2 inst_616 ( .SI(net_8379), .Q(net_8379), .SE(net_3969), .D(net_3937), .CK(net_10760) );
CLKBUF_X2 inst_10683 ( .A(net_10530), .Z(net_10531) );
CLKBUF_X2 inst_18293 ( .A(net_18140), .Z(net_18141) );
INV_X4 inst_5381 ( .ZN(net_1479), .A(net_1113) );
SDFF_X2 inst_1784 ( .D(net_7286), .SI(net_6903), .Q(net_6903), .SE(net_6284), .CK(net_16208) );
CLKBUF_X2 inst_18670 ( .A(net_18517), .Z(net_18518) );
AOI22_X2 inst_8040 ( .B1(net_7932), .A1(net_7830), .B2(net_6103), .A2(net_4398), .ZN(net_4099) );
CLKBUF_X2 inst_16402 ( .A(net_16249), .Z(net_16250) );
SDFFS_X2 inst_2071 ( .SI(net_7385), .SE(net_2795), .Q(net_174), .D(net_174), .CK(net_17498), .SN(x6501) );
CLKBUF_X2 inst_14921 ( .A(net_12320), .Z(net_14769) );
SDFF_X2 inst_1427 ( .SI(net_7287), .Q(net_7064), .D(net_7064), .SE(net_6280), .CK(net_18798) );
CLKBUF_X2 inst_10421 ( .A(net_9172), .Z(net_10269) );
AND2_X2 inst_9183 ( .A2(net_6093), .ZN(net_5988), .A1(net_2071) );
DFFR_X2 inst_7259 ( .QN(net_7400), .D(net_1978), .CK(net_17864), .RN(x6501) );
CLKBUF_X2 inst_10056 ( .A(net_9903), .Z(net_9904) );
CLKBUF_X2 inst_17346 ( .A(net_17193), .Z(net_17194) );
NAND2_X2 inst_4662 ( .ZN(net_2496), .A1(net_2230), .A2(net_2229) );
CLKBUF_X2 inst_14296 ( .A(net_14143), .Z(net_14144) );
XOR2_X1 inst_87 ( .A(net_2986), .Z(net_1931), .B(x3561) );
CLKBUF_X2 inst_17704 ( .A(net_17551), .Z(net_17552) );
CLKBUF_X2 inst_16172 ( .A(net_11650), .Z(net_16020) );
OAI22_X2 inst_2918 ( .ZN(net_3578), .A2(net_3212), .B1(net_3190), .B2(net_2203), .A1(net_1601) );
CLKBUF_X2 inst_10036 ( .A(net_9883), .Z(net_9884) );
SDFFR_X1 inst_2721 ( .SI(net_9031), .Q(net_9031), .D(net_7460), .SE(net_3208), .CK(net_10673), .RN(x6501) );
CLKBUF_X2 inst_9576 ( .A(net_9423), .Z(net_9424) );
OAI21_X2 inst_3074 ( .ZN(net_3904), .A(net_3902), .B2(net_3901), .B1(net_1156) );
SDFF_X2 inst_800 ( .SI(net_8339), .Q(net_8339), .D(net_3965), .SE(net_3880), .CK(net_10706) );
INV_X4 inst_5281 ( .ZN(net_1883), .A(net_1635) );
XOR2_X2 inst_10 ( .B(net_1794), .A(net_1790), .Z(net_1680) );
CLKBUF_X2 inst_9925 ( .A(net_9772), .Z(net_9773) );
AOI22_X2 inst_7770 ( .B1(net_6997), .A1(net_6957), .A2(net_5443), .B2(net_5442), .ZN(net_5323) );
NAND2_X2 inst_4337 ( .A1(net_7063), .A2(net_5162), .ZN(net_5120) );
CLKBUF_X2 inst_15550 ( .A(net_15397), .Z(net_15398) );
CLKBUF_X2 inst_10475 ( .A(net_10322), .Z(net_10323) );
AOI22_X2 inst_7981 ( .B1(net_7925), .A1(net_7823), .B2(net_6103), .A2(net_4398), .ZN(net_4150) );
CLKBUF_X2 inst_13555 ( .A(net_10605), .Z(net_13403) );
INV_X4 inst_5459 ( .ZN(net_881), .A(net_769) );
CLKBUF_X2 inst_13186 ( .A(net_9489), .Z(net_13034) );
CLKBUF_X2 inst_9867 ( .A(net_9225), .Z(net_9715) );
CLKBUF_X2 inst_18281 ( .A(net_15362), .Z(net_18129) );
CLKBUF_X2 inst_10090 ( .A(net_9791), .Z(net_9938) );
CLKBUF_X2 inst_16623 ( .A(net_12312), .Z(net_16471) );
CLKBUF_X2 inst_11961 ( .A(net_11808), .Z(net_11809) );
CLKBUF_X2 inst_16443 ( .A(net_10291), .Z(net_16291) );
CLKBUF_X2 inst_18368 ( .A(net_18215), .Z(net_18216) );
HA_X1 inst_6700 ( .CO(net_6105), .A(net_6078), .S(net_2463), .B(net_2462) );
CLKBUF_X2 inst_14462 ( .A(net_14309), .Z(net_14310) );
CLKBUF_X2 inst_16078 ( .A(net_15422), .Z(net_15926) );
NAND2_X2 inst_4731 ( .ZN(net_2708), .A2(net_1586), .A1(net_1226) );
SDFF_X2 inst_1276 ( .Q(net_7808), .D(net_7808), .SE(net_2730), .SI(net_2705), .CK(net_15853) );
XNOR2_X2 inst_256 ( .A(net_2668), .B(net_2512), .ZN(net_1193) );
INV_X2 inst_6205 ( .ZN(net_5505), .A(net_5409) );
SDFF_X2 inst_1902 ( .D(net_7297), .SI(net_7034), .Q(net_7034), .SE(net_6277), .CK(net_15403) );
AND2_X2 inst_9180 ( .ZN(net_2229), .A1(net_2139), .A2(net_2138) );
CLKBUF_X2 inst_16518 ( .A(net_16365), .Z(net_16366) );
AOI222_X1 inst_8626 ( .A2(net_8218), .C2(net_6117), .A1(net_4800), .B2(net_4799), .ZN(net_4798), .B1(net_3145), .C1(net_2205) );
CLKBUF_X2 inst_9635 ( .A(net_9482), .Z(net_9483) );
INV_X8 inst_5052 ( .ZN(net_6252), .A(net_3382) );
CLKBUF_X2 inst_16874 ( .A(net_16721), .Z(net_16722) );
INV_X4 inst_6038 ( .A(net_7361), .ZN(net_1750) );
CLKBUF_X2 inst_13791 ( .A(net_13638), .Z(net_13639) );
NAND3_X2 inst_3978 ( .A2(net_6117), .ZN(net_2078), .A1(net_2077), .A3(net_1769) );
INV_X4 inst_6106 ( .A(net_6366), .ZN(net_966) );
CLKBUF_X2 inst_11264 ( .A(net_11111), .Z(net_11112) );
CLKBUF_X2 inst_9354 ( .A(net_9201), .Z(net_9202) );
CLKBUF_X2 inst_10042 ( .A(net_9889), .Z(net_9890) );
CLKBUF_X2 inst_10214 ( .A(net_9081), .Z(net_10062) );
SDFFS_X2 inst_2078 ( .SI(net_7389), .SE(net_2795), .Q(net_178), .D(net_178), .CK(net_14664), .SN(x6501) );
AND2_X2 inst_9161 ( .ZN(net_2805), .A2(net_2804), .A1(net_2540) );
INV_X2 inst_6555 ( .A(net_8952), .ZN(net_500) );
CLKBUF_X2 inst_18773 ( .A(net_10541), .Z(net_18621) );
CLKBUF_X2 inst_17422 ( .A(net_10518), .Z(net_17270) );
SDFF_X2 inst_1462 ( .SI(net_7285), .Q(net_7142), .D(net_7142), .SE(net_6279), .CK(net_16215) );
AOI22_X2 inst_8509 ( .B1(net_6748), .A1(net_6715), .B2(net_6202), .A2(net_3520), .ZN(net_3431) );
SDFFR_X2 inst_2273 ( .D(net_7383), .SE(net_2797), .SI(net_192), .Q(net_192), .CK(net_14967), .RN(x6501) );
AND2_X4 inst_9138 ( .ZN(net_1385), .A2(net_795), .A1(net_178) );
INV_X2 inst_6391 ( .ZN(net_1257), .A(net_1256) );
CLKBUF_X2 inst_13944 ( .A(net_13791), .Z(net_13792) );
SDFF_X2 inst_2003 ( .SI(net_7784), .Q(net_7784), .D(net_2574), .SE(net_2459), .CK(net_16019) );
CLKBUF_X2 inst_15954 ( .A(net_15801), .Z(net_15802) );
INV_X4 inst_6100 ( .A(net_7371), .ZN(net_1121) );
INV_X4 inst_6084 ( .A(net_5974), .ZN(x3451) );
INV_X4 inst_5430 ( .ZN(net_2666), .A(net_832) );
INV_X4 inst_5119 ( .A(net_8228), .ZN(net_4628) );
MUX2_X2 inst_4963 ( .A(net_7387), .S(net_2370), .Z(net_2360), .B(net_787) );
SDFFR_X1 inst_2787 ( .D(net_7394), .Q(net_7291), .SI(net_1958), .SE(net_1327), .CK(net_15366), .RN(x6501) );
INV_X4 inst_5612 ( .A(net_6822), .ZN(net_1221) );
CLKBUF_X2 inst_13638 ( .A(net_13485), .Z(net_13486) );
CLKBUF_X2 inst_12455 ( .A(net_12302), .Z(net_12303) );
CLKBUF_X2 inst_9386 ( .A(net_9233), .Z(net_9234) );
CLKBUF_X2 inst_11074 ( .A(net_10921), .Z(net_10922) );
SDFFR_X2 inst_2599 ( .D(net_7376), .QN(net_7236), .SI(net_1866), .SE(net_1379), .CK(net_14647), .RN(x6501) );
CLKBUF_X2 inst_16062 ( .A(net_15909), .Z(net_15910) );
INV_X2 inst_6254 ( .ZN(net_4829), .A(net_4718) );
CLKBUF_X2 inst_18286 ( .A(net_11665), .Z(net_18134) );
NAND3_X2 inst_3971 ( .ZN(net_2385), .A1(net_2315), .A2(net_2164), .A3(net_2069) );
CLKBUF_X2 inst_11573 ( .A(net_10481), .Z(net_11421) );
CLKBUF_X2 inst_9858 ( .A(net_9705), .Z(net_9706) );
CLKBUF_X2 inst_18772 ( .A(net_18619), .Z(net_18620) );
CLKBUF_X2 inst_13596 ( .A(net_13443), .Z(net_13444) );
CLKBUF_X2 inst_18013 ( .A(net_16126), .Z(net_17861) );
SDFF_X2 inst_1123 ( .D(net_7329), .SI(net_6571), .Q(net_6571), .SE(net_3070), .CK(net_9511) );
CLKBUF_X2 inst_18028 ( .A(net_10515), .Z(net_17876) );
AOI221_X2 inst_8747 ( .ZN(net_5652), .A(net_5529), .B2(net_5520), .C2(net_4965), .B1(net_282), .C1(net_273) );
CLKBUF_X2 inst_13383 ( .A(net_12884), .Z(net_13231) );
CLKBUF_X2 inst_17256 ( .A(net_17103), .Z(net_17104) );
CLKBUF_X2 inst_11763 ( .A(net_11610), .Z(net_11611) );
DFFR_X2 inst_7169 ( .D(net_2579), .QN(net_342), .CK(net_11616), .RN(x6501) );
CLKBUF_X2 inst_16429 ( .A(net_11859), .Z(net_16277) );
AOI22_X2 inst_8061 ( .B1(net_8105), .A1(net_7765), .B2(net_6108), .A2(net_6096), .ZN(net_4081) );
SDFF_X2 inst_1628 ( .Q(net_8172), .D(net_8172), .SI(net_2710), .SE(net_2538), .CK(net_17130) );
DFF_X1 inst_6844 ( .Q(net_6434), .D(net_3603), .CK(net_17965) );
CLKBUF_X2 inst_17506 ( .A(net_17353), .Z(net_17354) );
CLKBUF_X2 inst_9640 ( .A(net_9374), .Z(net_9488) );
NAND2_X2 inst_4840 ( .A2(net_9009), .ZN(net_2429), .A1(net_557) );
XNOR2_X2 inst_225 ( .A(net_6363), .ZN(net_1364), .B(net_1363) );
CLKBUF_X2 inst_12530 ( .A(net_11125), .Z(net_12378) );
CLKBUF_X2 inst_14261 ( .A(net_14108), .Z(net_14109) );
CLKBUF_X2 inst_17832 ( .A(net_17679), .Z(net_17680) );
INV_X8 inst_5020 ( .ZN(net_5456), .A(net_4321) );
AND4_X4 inst_9030 ( .A2(net_7524), .ZN(net_1821), .A4(net_1705), .A3(net_1653), .A1(net_625) );
DFFR_X2 inst_7349 ( .Q(net_7318), .CK(net_11379), .D(x13115), .RN(x6501) );
CLKBUF_X2 inst_14808 ( .A(net_14445), .Z(net_14656) );
SDFF_X2 inst_508 ( .Q(net_8852), .D(net_8852), .SI(net_3961), .SE(net_3936), .CK(net_13204) );
NAND2_X2 inst_4888 ( .A2(net_7389), .ZN(net_708), .A1(net_178) );
AOI22_X2 inst_8150 ( .B1(net_8120), .A1(net_7882), .A2(net_6098), .B2(net_4190), .ZN(net_4002) );
CLKBUF_X2 inst_12611 ( .A(net_12458), .Z(net_12459) );
SDFF_X2 inst_590 ( .SI(net_8381), .Q(net_8381), .SE(net_3969), .D(net_3960), .CK(net_13126) );
SDFFR_X2 inst_2553 ( .QN(net_6360), .SE(net_2147), .D(net_2131), .SI(net_1956), .CK(net_17534), .RN(x6501) );
CLKBUF_X2 inst_18427 ( .A(net_18274), .Z(net_18275) );
CLKBUF_X2 inst_12209 ( .A(net_12056), .Z(net_12057) );
CLKBUF_X2 inst_12671 ( .A(net_12518), .Z(net_12519) );
CLKBUF_X2 inst_13051 ( .A(net_12898), .Z(net_12899) );
CLKBUF_X2 inst_13897 ( .A(net_13744), .Z(net_13745) );
NAND2_X2 inst_4531 ( .ZN(net_3382), .A2(net_3381), .A1(net_3378) );
SDFF_X2 inst_1105 ( .D(net_7335), .SI(net_6544), .Q(net_6544), .SE(net_3086), .CK(net_9755) );
SDFFR_X1 inst_2746 ( .SI(net_9040), .Q(net_9040), .D(net_7469), .SE(net_3208), .CK(net_12202), .RN(x6501) );
CLKBUF_X2 inst_14746 ( .A(net_13929), .Z(net_14594) );
CLKBUF_X2 inst_14387 ( .A(net_14234), .Z(net_14235) );
DFFS_X1 inst_6961 ( .D(net_1687), .CK(net_16328), .SN(x6501), .Q(x956) );
AOI22_X2 inst_8200 ( .B1(net_8829), .A1(net_8348), .A2(net_6265), .B2(net_6253), .ZN(net_3836) );
XNOR2_X2 inst_330 ( .B(net_7373), .A(net_6355), .ZN(net_819) );
CLKBUF_X2 inst_13345 ( .A(net_13192), .Z(net_13193) );
CLKBUF_X2 inst_13558 ( .A(net_13405), .Z(net_13406) );
NAND2_X2 inst_4305 ( .A1(net_7134), .A2(net_5166), .ZN(net_5152) );
CLKBUF_X2 inst_12101 ( .A(net_9215), .Z(net_11949) );
CLKBUF_X2 inst_13546 ( .A(net_13393), .Z(net_13394) );
AOI221_X2 inst_8786 ( .B1(net_7200), .C2(net_6130), .B2(net_5655), .ZN(net_5037), .A(net_4772), .C1(net_1298) );
NOR2_X2 inst_3566 ( .A1(net_6752), .ZN(net_2905), .A2(net_1465) );
CLKBUF_X2 inst_13864 ( .A(net_13028), .Z(net_13712) );
CLKBUF_X2 inst_11803 ( .A(net_11466), .Z(net_11651) );
CLKBUF_X2 inst_15455 ( .A(net_15302), .Z(net_15303) );
CLKBUF_X2 inst_16108 ( .A(net_15955), .Z(net_15956) );
SDFF_X2 inst_1232 ( .Q(net_7826), .D(net_7826), .SE(net_2730), .SI(net_2718), .CK(net_15634) );
CLKBUF_X2 inst_14431 ( .A(net_14278), .Z(net_14279) );
CLKBUF_X2 inst_16562 ( .A(net_16409), .Z(net_16410) );
CLKBUF_X2 inst_18968 ( .A(net_12588), .Z(net_18816) );
SDFF_X2 inst_758 ( .Q(net_8799), .D(net_8799), .SI(net_3956), .SE(net_3879), .CK(net_10902) );
CLKBUF_X2 inst_17915 ( .A(net_17762), .Z(net_17763) );
SDFFR_X2 inst_2146 ( .Q(net_8891), .D(net_8891), .SE(net_3901), .SI(net_1408), .CK(net_13510), .RN(x6501) );
CLKBUF_X2 inst_13332 ( .A(net_13179), .Z(net_13180) );
AOI22_X2 inst_8543 ( .B1(net_6594), .A1(net_6561), .A2(net_6257), .B2(net_6110), .ZN(net_3397) );
NOR2_X2 inst_3437 ( .A2(net_3093), .ZN(net_3067), .A1(net_2302) );
CLKBUF_X2 inst_13425 ( .A(net_13272), .Z(net_13273) );
DFF_X1 inst_6813 ( .Q(net_8218), .D(net_4454), .CK(net_14461) );
CLKBUF_X2 inst_17777 ( .A(net_17624), .Z(net_17625) );
INV_X4 inst_5764 ( .A(net_9007), .ZN(net_2680) );
DFFR_X1 inst_7442 ( .QN(net_8921), .D(net_4762), .CK(net_13971), .RN(x6501) );
SDFF_X2 inst_1953 ( .D(net_7271), .SI(net_6888), .Q(net_6888), .SE(net_6284), .CK(net_14077) );
NAND2_X2 inst_4570 ( .A2(net_6200), .A1(net_6106), .ZN(net_3059) );
OAI21_X2 inst_3016 ( .ZN(net_5046), .B2(net_5044), .A(net_4893), .B1(net_1485) );
SDFF_X2 inst_1958 ( .D(net_7270), .SI(net_6887), .Q(net_6887), .SE(net_6284), .CK(net_14318) );
CLKBUF_X2 inst_14050 ( .A(net_13897), .Z(net_13898) );
CLKBUF_X2 inst_18639 ( .A(net_11333), .Z(net_18487) );
DFFS_X2 inst_6885 ( .Q(net_8256), .D(net_3179), .CK(net_18469), .SN(x6501) );
NOR4_X2 inst_3240 ( .A4(net_7367), .A3(net_7366), .ZN(net_1835), .A2(net_1625), .A1(net_893) );
CLKBUF_X2 inst_9403 ( .A(net_9250), .Z(net_9251) );
CLKBUF_X2 inst_17201 ( .A(net_17048), .Z(net_17049) );
CLKBUF_X2 inst_16950 ( .A(net_9768), .Z(net_16798) );
CLKBUF_X2 inst_19022 ( .A(net_18869), .Z(net_18870) );
XNOR2_X2 inst_111 ( .A(net_6267), .ZN(net_4682), .B(net_4355) );
CLKBUF_X2 inst_13196 ( .A(net_13043), .Z(net_13044) );
SDFF_X2 inst_1723 ( .SI(net_7268), .Q(net_7045), .D(net_7045), .SE(net_6280), .CK(net_14360) );
NOR3_X2 inst_3278 ( .ZN(net_2789), .A1(net_2400), .A3(net_2398), .A2(net_2397) );
CLKBUF_X2 inst_11425 ( .A(net_11272), .Z(net_11273) );
INV_X4 inst_5145 ( .ZN(net_6055), .A(net_3304) );
CLKBUF_X2 inst_11296 ( .A(net_11143), .Z(net_11144) );
CLKBUF_X2 inst_16703 ( .A(net_16550), .Z(net_16551) );
CLKBUF_X2 inst_13407 ( .A(net_11512), .Z(net_13255) );
CLKBUF_X2 inst_17906 ( .A(net_13433), .Z(net_17754) );
SDFF_X2 inst_978 ( .SI(net_7342), .Q(net_6749), .D(net_6749), .SE(net_3124), .CK(net_11688) );
CLKBUF_X2 inst_14757 ( .A(net_14604), .Z(net_14605) );
OAI221_X2 inst_2955 ( .ZN(net_4923), .B1(net_4922), .C2(net_4774), .B2(net_4530), .A(net_2889), .C1(net_1520) );
CLKBUF_X2 inst_13506 ( .A(net_13041), .Z(net_13354) );
NAND3_X2 inst_3926 ( .ZN(net_5612), .A1(net_5541), .A3(net_5475), .A2(net_5287) );
DFFR_X2 inst_7293 ( .D(net_7618), .QN(net_7617), .CK(net_17994), .RN(x6501) );
CLKBUF_X2 inst_16515 ( .A(net_9274), .Z(net_16363) );
CLKBUF_X2 inst_13160 ( .A(net_9660), .Z(net_13008) );
CLKBUF_X2 inst_17765 ( .A(net_15275), .Z(net_17613) );
CLKBUF_X2 inst_9745 ( .A(net_9592), .Z(net_9593) );
CLKBUF_X2 inst_18295 ( .A(net_18142), .Z(net_18143) );
CLKBUF_X2 inst_19030 ( .A(net_15046), .Z(net_18878) );
SDFF_X2 inst_495 ( .SI(net_8620), .Q(net_8620), .SE(net_3984), .D(net_3941), .CK(net_13430) );
CLKBUF_X2 inst_14366 ( .A(net_14116), .Z(net_14214) );
CLKBUF_X2 inst_15041 ( .A(net_14888), .Z(net_14889) );
INV_X2 inst_6437 ( .A(net_1568), .ZN(net_657) );
SDFF_X2 inst_1864 ( .D(net_7298), .SI(net_6955), .Q(net_6955), .SE(net_6281), .CK(net_18182) );
CLKBUF_X2 inst_9632 ( .A(net_9479), .Z(net_9480) );
NOR4_X2 inst_3224 ( .ZN(net_2384), .A1(net_2118), .A2(net_1746), .A4(net_987), .A3(net_979) );
CLKBUF_X2 inst_16626 ( .A(net_14056), .Z(net_16474) );
CLKBUF_X2 inst_10887 ( .A(net_10734), .Z(net_10735) );
CLKBUF_X2 inst_18534 ( .A(net_18381), .Z(net_18382) );
AOI22_X2 inst_7917 ( .A1(net_8993), .A2(net_5456), .B2(net_5260), .ZN(net_4466), .B1(net_4465) );
CLKBUF_X2 inst_12616 ( .A(net_12463), .Z(net_12464) );
CLKBUF_X2 inst_15826 ( .A(net_15673), .Z(net_15674) );
CLKBUF_X2 inst_16852 ( .A(net_16699), .Z(net_16700) );
CLKBUF_X2 inst_13305 ( .A(net_13152), .Z(net_13153) );
DFFR_X2 inst_7286 ( .QN(net_6345), .D(net_1610), .CK(net_15182), .RN(x6501) );
CLKBUF_X2 inst_12644 ( .A(net_12491), .Z(net_12492) );
AOI21_X2 inst_8914 ( .B2(net_5871), .ZN(net_5724), .A(net_5721), .B1(x480) );
CLKBUF_X2 inst_18150 ( .A(net_17997), .Z(net_17998) );
OR2_X2 inst_2893 ( .A1(net_7303), .ZN(net_1685), .A2(net_1631) );
CLKBUF_X2 inst_9497 ( .A(net_9344), .Z(net_9345) );
DFF_X1 inst_6727 ( .Q(net_6773), .D(net_5642), .CK(net_9221) );
CLKBUF_X2 inst_12447 ( .A(net_12294), .Z(net_12295) );
AOI22_X2 inst_7937 ( .B1(net_8020), .A1(net_7986), .B2(net_6102), .A2(net_6097), .ZN(net_4187) );
INV_X2 inst_6347 ( .A(net_2945), .ZN(net_2518) );
SDFF_X2 inst_1453 ( .SI(net_7271), .Q(net_7088), .D(net_7088), .SE(net_6278), .CK(net_16848) );
CLKBUF_X2 inst_12466 ( .A(net_12313), .Z(net_12314) );
AOI21_X2 inst_8871 ( .B2(net_6254), .ZN(net_5936), .A(net_5934), .B1(x1070) );
CLKBUF_X2 inst_17961 ( .A(net_17808), .Z(net_17809) );
OAI21_X2 inst_3007 ( .B2(net_5755), .ZN(net_5743), .A(net_5740), .B1(net_563) );
CLKBUF_X2 inst_18344 ( .A(net_15414), .Z(net_18192) );
CLKBUF_X2 inst_15081 ( .A(net_14928), .Z(net_14929) );
NAND2_X2 inst_4185 ( .ZN(net_5317), .A1(net_5071), .A2(net_5070) );
INV_X2 inst_6358 ( .ZN(net_2190), .A(net_2100) );
NOR2_X2 inst_3512 ( .A2(net_4391), .ZN(net_1805), .A1(net_1658) );
CLKBUF_X2 inst_11018 ( .A(net_10865), .Z(net_10866) );
CLKBUF_X2 inst_11485 ( .A(net_11332), .Z(net_11333) );
CLKBUF_X2 inst_10738 ( .A(net_10585), .Z(net_10586) );
INV_X4 inst_5632 ( .A(net_6314), .ZN(net_2726) );
CLKBUF_X2 inst_14839 ( .A(net_14686), .Z(net_14687) );
SDFF_X2 inst_1206 ( .Q(net_7825), .D(net_7825), .SE(net_2730), .SI(net_2722), .CK(net_17725) );
CLKBUF_X2 inst_15778 ( .A(net_15625), .Z(net_15626) );
CLKBUF_X2 inst_15270 ( .A(net_15117), .Z(net_15118) );
DFF_X1 inst_6773 ( .Q(net_7552), .D(net_4599), .CK(net_10483) );
CLKBUF_X2 inst_15485 ( .A(net_15332), .Z(net_15333) );
DFFR_X2 inst_7075 ( .QN(net_8296), .D(net_3972), .CK(net_11244), .RN(x6501) );
CLKBUF_X2 inst_10328 ( .A(net_10175), .Z(net_10176) );
NOR2_X2 inst_3466 ( .A1(net_6121), .ZN(net_4800), .A2(net_2474) );
AOI22_X2 inst_8106 ( .A1(net_7975), .B1(net_7805), .A2(net_6092), .B2(net_6091), .ZN(net_4041) );
AOI22_X2 inst_8358 ( .B1(net_8591), .A1(net_8480), .A2(net_6263), .B2(net_6262), .ZN(net_3690) );
CLKBUF_X2 inst_13907 ( .A(net_13754), .Z(net_13755) );
NAND2_X2 inst_4800 ( .ZN(net_1632), .A2(net_1376), .A1(net_1267) );
NAND2_X2 inst_4394 ( .A1(net_7044), .A2(net_5162), .ZN(net_5063) );
CLKBUF_X2 inst_15684 ( .A(net_15531), .Z(net_15532) );
CLKBUF_X2 inst_11303 ( .A(net_9269), .Z(net_11151) );
CLKBUF_X2 inst_12631 ( .A(net_12478), .Z(net_12479) );
CLKBUF_X2 inst_13086 ( .A(net_10631), .Z(net_12934) );
SDFF_X2 inst_1487 ( .SI(net_7284), .Q(net_7061), .D(net_7061), .SE(net_6280), .CK(net_16212) );
AOI22_X2 inst_7807 ( .A2(net_8218), .B2(net_6144), .ZN(net_4766), .A1(net_4764), .B1(net_4528) );
DFFR_X2 inst_7246 ( .QN(net_7403), .D(net_2053), .CK(net_17870), .RN(x6501) );
SDFF_X2 inst_1933 ( .SI(net_8063), .Q(net_8063), .D(net_2722), .SE(net_2508), .CK(net_18749) );
CLKBUF_X2 inst_13169 ( .A(net_13016), .Z(net_13017) );
DFFR_X1 inst_7511 ( .Q(net_6338), .D(net_1505), .CK(net_14844), .RN(x6501) );
CLKBUF_X2 inst_18996 ( .A(net_14745), .Z(net_18844) );
CLKBUF_X2 inst_12025 ( .A(net_11872), .Z(net_11873) );
NAND2_X2 inst_4320 ( .A1(net_7139), .A2(net_5166), .ZN(net_5137) );
CLKBUF_X2 inst_16120 ( .A(net_14640), .Z(net_15968) );
CLKBUF_X2 inst_16031 ( .A(net_15878), .Z(net_15879) );
DFFR_X1 inst_7572 ( .Q(net_7643), .D(net_7634), .CK(net_15697), .RN(x6501) );
INV_X2 inst_6313 ( .A(net_3552), .ZN(net_3548) );
CLKBUF_X2 inst_16810 ( .A(net_16657), .Z(net_16658) );
CLKBUF_X2 inst_18101 ( .A(net_17948), .Z(net_17949) );
CLKBUF_X2 inst_15516 ( .A(net_15215), .Z(net_15364) );
CLKBUF_X2 inst_14228 ( .A(net_11128), .Z(net_14076) );
CLKBUF_X2 inst_14316 ( .A(net_14163), .Z(net_14164) );
CLKBUF_X2 inst_14182 ( .A(net_13150), .Z(net_14030) );
NAND2_X2 inst_4771 ( .A1(net_7618), .A2(net_7617), .ZN(net_2777) );
CLKBUF_X2 inst_16986 ( .A(net_16833), .Z(net_16834) );
CLKBUF_X2 inst_16375 ( .A(net_13106), .Z(net_16223) );
NAND2_X2 inst_4669 ( .ZN(net_2398), .A2(net_2162), .A1(net_1598) );
CLKBUF_X2 inst_15091 ( .A(net_12208), .Z(net_14939) );
CLKBUF_X2 inst_15476 ( .A(net_15323), .Z(net_15324) );
AOI22_X2 inst_8016 ( .B1(net_8099), .A1(net_7759), .B2(net_6108), .A2(net_6096), .ZN(net_4120) );
AOI221_X4 inst_8707 ( .C1(net_8197), .B1(net_7687), .C2(net_6099), .ZN(net_6037), .B2(net_4399), .A(net_4302) );
CLKBUF_X2 inst_13204 ( .A(net_11873), .Z(net_13052) );
CLKBUF_X2 inst_15191 ( .A(net_12457), .Z(net_15039) );
CLKBUF_X2 inst_12230 ( .A(net_10247), .Z(net_12078) );
CLKBUF_X2 inst_15650 ( .A(net_15497), .Z(net_15498) );
SDFF_X2 inst_1017 ( .SI(net_7331), .Q(net_6672), .D(net_6672), .SE(net_3126), .CK(net_9432) );
CLKBUF_X2 inst_13802 ( .A(net_10325), .Z(net_13650) );
XNOR2_X2 inst_281 ( .ZN(net_1022), .A(net_1021), .B(net_1020) );
INV_X2 inst_6336 ( .ZN(net_2884), .A(net_2837) );
CLKBUF_X2 inst_10306 ( .A(net_9553), .Z(net_10154) );
DFFR_X2 inst_7062 ( .QN(net_7174), .D(net_4313), .CK(net_13602), .RN(x6501) );
SDFF_X2 inst_1836 ( .D(net_7274), .SI(net_6891), .Q(net_6891), .SE(net_6284), .CK(net_14114) );
CLKBUF_X2 inst_18103 ( .A(net_17950), .Z(net_17951) );
DFFR_X2 inst_7005 ( .D(net_5878), .CK(net_9226), .RN(x6501), .Q(x2261) );
NAND2_X2 inst_4274 ( .A1(net_7039), .A2(net_5249), .ZN(net_5186) );
NAND2_X2 inst_4250 ( .A1(net_7028), .A2(net_5249), .ZN(net_5210) );
SDFFR_X2 inst_2170 ( .QN(net_7567), .D(net_3947), .SE(net_3144), .SI(net_3131), .CK(net_13219), .RN(x6501) );
DFFR_X1 inst_7414 ( .D(net_5727), .CK(net_13823), .RN(x6501), .Q(x27) );
CLKBUF_X2 inst_13322 ( .A(net_9691), .Z(net_13170) );
CLKBUF_X2 inst_15490 ( .A(net_15337), .Z(net_15338) );
OAI22_X2 inst_2946 ( .A1(net_7526), .B2(net_7524), .A2(net_6325), .ZN(net_1702), .B1(net_1700) );
CLKBUF_X2 inst_9940 ( .A(net_9787), .Z(net_9788) );
CLKBUF_X2 inst_14149 ( .A(net_13996), .Z(net_13997) );
CLKBUF_X2 inst_16415 ( .A(net_16262), .Z(net_16263) );
CLKBUF_X2 inst_15234 ( .A(net_13547), .Z(net_15082) );
CLKBUF_X2 inst_13827 ( .A(net_13674), .Z(net_13675) );
CLKBUF_X2 inst_10828 ( .A(net_10675), .Z(net_10676) );
CLKBUF_X2 inst_18932 ( .A(net_18779), .Z(net_18780) );
OAI211_X2 inst_3211 ( .C2(net_6820), .ZN(net_2283), .B(net_2282), .C1(net_2015), .A(net_1393) );
CLKBUF_X2 inst_10364 ( .A(net_9206), .Z(net_10212) );
CLKBUF_X2 inst_12702 ( .A(net_12549), .Z(net_12550) );
DFFR_X2 inst_7270 ( .QN(net_7231), .D(net_1987), .CK(net_14776), .RN(x6501) );
CLKBUF_X2 inst_10906 ( .A(net_10753), .Z(net_10754) );
CLKBUF_X2 inst_14803 ( .A(net_14650), .Z(net_14651) );
CLKBUF_X2 inst_18415 ( .A(net_18262), .Z(net_18263) );
SDFFR_X2 inst_2386 ( .SE(net_2260), .Q(net_373), .D(net_373), .CK(net_11454), .RN(x6501), .SI(x1575) );
CLKBUF_X2 inst_13846 ( .A(net_13693), .Z(net_13694) );
NAND2_X2 inst_4103 ( .ZN(net_5429), .A1(net_5241), .A2(net_5013) );
SDFF_X2 inst_1267 ( .Q(net_8086), .D(net_8086), .SE(net_2707), .SI(net_2702), .CK(net_18895) );
SDFF_X2 inst_1507 ( .SI(net_7868), .Q(net_7868), .D(net_2715), .SE(net_2558), .CK(net_16828) );
CLKBUF_X2 inst_15276 ( .A(net_15123), .Z(net_15124) );
CLKBUF_X2 inst_19116 ( .A(net_9700), .Z(net_18964) );
CLKBUF_X2 inst_19091 ( .A(net_18938), .Z(net_18939) );
DFFR_X2 inst_7301 ( .D(net_6419), .Q(net_6414), .CK(net_18708), .RN(x6501) );
DFFR_X2 inst_7260 ( .QN(net_7235), .D(net_1981), .CK(net_14784), .RN(x6501) );
NAND4_X2 inst_3786 ( .ZN(net_4235), .A1(net_3663), .A2(net_3662), .A3(net_3661), .A4(net_3660) );
CLKBUF_X2 inst_14960 ( .A(net_14807), .Z(net_14808) );
DFFR_X1 inst_7367 ( .D(net_5938), .CK(net_11987), .RN(x6501), .Q(x1070) );
NOR2_X2 inst_3404 ( .A2(net_6145), .ZN(net_3877), .A1(net_3323) );
AOI22_X2 inst_7878 ( .B2(net_4881), .A2(net_4809), .ZN(net_4561), .A1(net_340), .B1(net_233) );
INV_X4 inst_5351 ( .A(net_2019), .ZN(net_1631) );
SDFF_X2 inst_542 ( .Q(net_8686), .D(net_8686), .SI(net_3974), .SE(net_3935), .CK(net_10166) );
XNOR2_X2 inst_128 ( .B(net_6318), .ZN(net_2858), .A(net_2536) );
CLKBUF_X2 inst_13589 ( .A(net_13436), .Z(net_13437) );
CLKBUF_X2 inst_18946 ( .A(net_18793), .Z(net_18794) );
CLKBUF_X2 inst_14172 ( .A(net_14019), .Z(net_14020) );
CLKBUF_X2 inst_14322 ( .A(net_14169), .Z(net_14170) );
CLKBUF_X2 inst_13100 ( .A(net_12947), .Z(net_12948) );
CLKBUF_X2 inst_13222 ( .A(net_13069), .Z(net_13070) );
CLKBUF_X2 inst_15252 ( .A(net_15099), .Z(net_15100) );
NAND3_X2 inst_4000 ( .ZN(net_4408), .A1(net_4322), .A3(net_1521), .A2(net_1149) );
CLKBUF_X2 inst_13625 ( .A(net_13472), .Z(net_13473) );
NOR4_X2 inst_3218 ( .ZN(net_5468), .A2(net_4838), .A1(net_4822), .A4(net_4775), .A3(net_2938) );
DFFS_X2 inst_6904 ( .QN(net_6819), .D(net_2016), .CK(net_18700), .SN(x6501) );
CLKBUF_X2 inst_9345 ( .A(net_9192), .Z(net_9193) );
AOI22_X2 inst_8137 ( .B1(net_7914), .A1(net_7812), .B2(net_6103), .A2(net_4398), .ZN(net_4013) );
INV_X4 inst_5723 ( .A(net_8933), .ZN(net_2598) );
OAI221_X2 inst_2958 ( .C2(net_8243), .B1(net_7586), .B2(net_4971), .C1(net_4928), .ZN(net_4845), .A(net_3389) );
XOR2_X2 inst_24 ( .A(net_6140), .B(net_4617), .Z(net_1365) );
SDFF_X2 inst_1209 ( .Q(net_7972), .D(net_7972), .SE(net_2755), .SI(net_2704), .CK(net_17040) );
CLKBUF_X2 inst_16832 ( .A(net_16679), .Z(net_16680) );
AOI22_X2 inst_8190 ( .B1(net_8680), .A1(net_8643), .B2(net_6109), .A2(net_3857), .ZN(net_3843) );
SDFF_X2 inst_1611 ( .Q(net_8118), .D(net_8118), .SI(net_2708), .SE(net_2541), .CK(net_18268) );
NAND2_X2 inst_4469 ( .ZN(net_4726), .A2(net_4725), .A1(net_4504) );
DFF_X1 inst_6779 ( .Q(net_7557), .D(net_4593), .CK(net_12757) );
CLKBUF_X2 inst_12764 ( .A(net_12611), .Z(net_12612) );
AOI221_X4 inst_8730 ( .B1(net_8846), .C1(net_8365), .C2(net_6265), .B2(net_6253), .ZN(net_4335), .A(net_4243) );
AOI22_X2 inst_8466 ( .B1(net_6672), .A1(net_6639), .A2(net_6213), .B2(net_6138), .ZN(net_3474) );
INV_X4 inst_5849 ( .A(net_7359), .ZN(net_1908) );
CLKBUF_X2 inst_17005 ( .A(net_16852), .Z(net_16853) );
SDFF_X2 inst_1663 ( .SI(net_7757), .Q(net_7757), .D(net_2722), .SE(net_2560), .CK(net_18772) );
SDFFR_X1 inst_2714 ( .Q(net_7633), .D(net_7633), .SE(net_3901), .SI(net_1157), .CK(net_13519), .RN(x6501) );
CLKBUF_X2 inst_13223 ( .A(net_10991), .Z(net_13071) );
DFFR_X2 inst_7099 ( .QN(net_6457), .D(net_3348), .CK(net_15100), .RN(x6501) );
CLKBUF_X2 inst_13036 ( .A(net_12883), .Z(net_12884) );
AOI22_X2 inst_7962 ( .B1(net_8058), .A1(net_7854), .B2(net_6107), .A2(net_4400), .ZN(net_4166) );
CLKBUF_X2 inst_15730 ( .A(net_15577), .Z(net_15578) );
CLKBUF_X2 inst_16029 ( .A(net_15876), .Z(net_15877) );
CLKBUF_X2 inst_15420 ( .A(net_15267), .Z(net_15268) );
CLKBUF_X2 inst_11285 ( .A(net_11132), .Z(net_11133) );
CLKBUF_X2 inst_10713 ( .A(net_10560), .Z(net_10561) );
CLKBUF_X2 inst_14928 ( .A(net_11766), .Z(net_14776) );
CLKBUF_X2 inst_15088 ( .A(net_14935), .Z(net_14936) );
CLKBUF_X2 inst_18929 ( .A(net_18776), .Z(net_18777) );
CLKBUF_X2 inst_16228 ( .A(net_16075), .Z(net_16076) );
INV_X4 inst_6021 ( .A(net_5978), .ZN(x3685) );
SDFF_X2 inst_820 ( .SI(net_8484), .Q(net_8484), .D(net_3980), .SE(net_3884), .CK(net_10695) );
XNOR2_X2 inst_157 ( .ZN(net_1940), .A(net_1680), .B(net_1640) );
SDFF_X2 inst_1441 ( .SI(net_7286), .Q(net_7103), .D(net_7103), .SE(net_6278), .CK(net_16222) );
OAI22_X2 inst_2929 ( .ZN(net_2523), .A2(net_2522), .A1(net_2312), .B2(net_2220), .B1(net_763) );
CLKBUF_X2 inst_12154 ( .A(net_10554), .Z(net_12002) );
NOR2_X2 inst_3443 ( .A2(net_3093), .ZN(net_3045), .A1(net_2745) );
INV_X4 inst_6159 ( .ZN(net_6207), .A(net_6206) );
NAND2_X2 inst_4287 ( .A1(net_6888), .A2(net_5247), .ZN(net_5173) );
CLKBUF_X2 inst_10986 ( .A(net_10833), .Z(net_10834) );
INV_X4 inst_5491 ( .ZN(net_834), .A(net_722) );
SDFFR_X2 inst_2177 ( .QN(net_7590), .D(net_3952), .SE(net_3144), .SI(net_714), .CK(net_10385), .RN(x6501) );
CLKBUF_X2 inst_16963 ( .A(net_9203), .Z(net_16811) );
CLKBUF_X2 inst_9588 ( .A(net_9435), .Z(net_9436) );
DFFR_X1 inst_7447 ( .QN(net_8922), .D(net_4761), .CK(net_14589), .RN(x6501) );
AOI22_X2 inst_8348 ( .B1(net_8590), .A1(net_8479), .A2(net_6263), .B2(net_6262), .ZN(net_3700) );
CLKBUF_X2 inst_17549 ( .A(net_11208), .Z(net_17397) );
NOR2_X2 inst_3410 ( .A2(net_6255), .ZN(net_3563), .A1(net_3304) );
INV_X4 inst_5339 ( .A(net_1479), .ZN(net_1311) );
CLKBUF_X2 inst_11506 ( .A(net_11353), .Z(net_11354) );
CLKBUF_X2 inst_13478 ( .A(net_13325), .Z(net_13326) );
CLKBUF_X2 inst_13216 ( .A(net_10531), .Z(net_13064) );
CLKBUF_X2 inst_17227 ( .A(net_17074), .Z(net_17075) );
XOR2_X2 inst_17 ( .Z(net_1422), .B(net_1421), .A(net_639) );
CLKBUF_X2 inst_10105 ( .A(net_9952), .Z(net_9953) );
AOI22_X2 inst_7838 ( .A1(net_7176), .A2(net_5655), .B2(net_5595), .ZN(net_4673), .B1(net_309) );
XNOR2_X2 inst_249 ( .A(net_2727), .B(net_2675), .ZN(net_1201) );
SDFFR_X2 inst_2234 ( .SI(net_9053), .Q(net_9053), .SE(net_2963), .D(net_1919), .CK(net_11126), .RN(x6501) );
CLKBUF_X2 inst_12407 ( .A(net_12254), .Z(net_12255) );
INV_X2 inst_6251 ( .ZN(net_4855), .A(net_4739) );
CLKBUF_X2 inst_18879 ( .A(net_18726), .Z(net_18727) );
CLKBUF_X2 inst_14509 ( .A(net_14356), .Z(net_14357) );
INV_X4 inst_5204 ( .ZN(net_5784), .A(net_5718) );
SDFF_X2 inst_1480 ( .SI(net_7267), .Q(net_7044), .D(net_7044), .SE(net_6280), .CK(net_16834) );
CLKBUF_X2 inst_18905 ( .A(net_18752), .Z(net_18753) );
CLKBUF_X2 inst_17461 ( .A(net_17308), .Z(net_17309) );
CLKBUF_X2 inst_10676 ( .A(net_10523), .Z(net_10524) );
CLKBUF_X2 inst_14121 ( .A(net_9301), .Z(net_13969) );
CLKBUF_X2 inst_15305 ( .A(net_15152), .Z(net_15153) );
CLKBUF_X2 inst_18856 ( .A(net_10228), .Z(net_18704) );
CLKBUF_X2 inst_17334 ( .A(net_17181), .Z(net_17182) );
CLKBUF_X2 inst_15708 ( .A(net_15555), .Z(net_15556) );
CLKBUF_X2 inst_17173 ( .A(net_17020), .Z(net_17021) );
CLKBUF_X2 inst_12359 ( .A(net_12206), .Z(net_12207) );
DFFR_X1 inst_7409 ( .D(net_5704), .CK(net_14038), .RN(x6501), .Q(x338) );
INV_X2 inst_6472 ( .A(net_7588), .ZN(net_3135) );
CLKBUF_X2 inst_10504 ( .A(net_10351), .Z(net_10352) );
CLKBUF_X2 inst_18450 ( .A(net_18297), .Z(net_18298) );
CLKBUF_X2 inst_16704 ( .A(net_16551), .Z(net_16552) );
SDFF_X2 inst_664 ( .Q(net_8438), .D(net_8438), .SI(net_3940), .SE(net_3934), .CK(net_13476) );
CLKBUF_X2 inst_11638 ( .A(net_9401), .Z(net_11486) );
CLKBUF_X2 inst_13977 ( .A(net_13824), .Z(net_13825) );
CLKBUF_X2 inst_10486 ( .A(net_10333), .Z(net_10334) );
CLKBUF_X2 inst_12485 ( .A(net_12196), .Z(net_12333) );
CLKBUF_X2 inst_14262 ( .A(net_14109), .Z(net_14110) );
CLKBUF_X2 inst_9911 ( .A(net_9758), .Z(net_9759) );
SDFF_X2 inst_1918 ( .D(net_7296), .SI(net_6913), .Q(net_6913), .SE(net_6284), .CK(net_15400) );
CLKBUF_X2 inst_9466 ( .A(net_9313), .Z(net_9314) );
CLKBUF_X2 inst_14500 ( .A(net_14347), .Z(net_14348) );
CLKBUF_X2 inst_17441 ( .A(net_12448), .Z(net_17289) );
CLKBUF_X2 inst_16590 ( .A(net_16187), .Z(net_16438) );
CLKBUF_X2 inst_15394 ( .A(net_15241), .Z(net_15242) );
NAND2_X2 inst_4064 ( .ZN(net_5875), .A2(net_5772), .A1(net_3234) );
NAND2_X2 inst_4427 ( .A1(net_6865), .A2(net_5016), .ZN(net_5000) );
CLKBUF_X2 inst_15806 ( .A(net_11003), .Z(net_15654) );
CLKBUF_X2 inst_12543 ( .A(net_12390), .Z(net_12391) );
NAND2_X2 inst_4635 ( .ZN(net_2835), .A1(net_2473), .A2(net_2325) );
NAND4_X2 inst_3839 ( .ZN(net_1967), .A3(net_1699), .A4(net_1251), .A2(net_1240), .A1(net_949) );
AOI22_X2 inst_7862 ( .B2(net_4881), .A2(net_4809), .ZN(net_4579), .A1(net_344), .B1(net_250) );
SDFFR_X2 inst_2368 ( .D(net_7366), .SE(net_2738), .SI(net_1916), .QN(net_262), .CK(net_13550), .RN(x6501) );
SDFFR_X1 inst_2735 ( .SI(net_5953), .Q(net_5953), .SE(net_3208), .D(net_3128), .CK(net_13511), .RN(x6501) );
OAI22_X2 inst_2934 ( .B1(net_8903), .ZN(net_2158), .A2(net_2157), .B2(net_2156), .A1(net_1923) );
SDFFR_X1 inst_2767 ( .Q(net_7295), .D(net_2073), .SI(net_1994), .SE(net_1327), .CK(net_18254), .RN(x6501) );
SDFF_X2 inst_1370 ( .SI(net_7282), .Q(net_7139), .D(net_7139), .SE(net_6279), .CK(net_14932) );
SDFFR_X2 inst_2512 ( .Q(net_7560), .D(net_7560), .SI(net_2760), .SE(net_2182), .CK(net_17802), .RN(x6501) );
CLKBUF_X2 inst_15805 ( .A(net_15652), .Z(net_15653) );
CLKBUF_X2 inst_12093 ( .A(net_11940), .Z(net_11941) );
CLKBUF_X2 inst_11948 ( .A(net_11795), .Z(net_11796) );
CLKBUF_X2 inst_17587 ( .A(net_17434), .Z(net_17435) );
CLKBUF_X2 inst_11447 ( .A(net_11294), .Z(net_11295) );
CLKBUF_X2 inst_18884 ( .A(net_18731), .Z(net_18732) );
CLKBUF_X2 inst_12568 ( .A(net_12415), .Z(net_12416) );
NAND2_X2 inst_4124 ( .ZN(net_5401), .A1(net_5227), .A2(net_5006) );
CLKBUF_X2 inst_13078 ( .A(net_12925), .Z(net_12926) );
CLKBUF_X2 inst_15886 ( .A(net_15580), .Z(net_15734) );
CLKBUF_X2 inst_14740 ( .A(net_14587), .Z(net_14588) );
CLKBUF_X2 inst_17648 ( .A(net_17495), .Z(net_17496) );
CLKBUF_X2 inst_15837 ( .A(net_15684), .Z(net_15685) );
INV_X4 inst_5672 ( .A(net_6288), .ZN(net_2728) );
CLKBUF_X2 inst_17987 ( .A(net_17834), .Z(net_17835) );
CLKBUF_X2 inst_10273 ( .A(net_10120), .Z(net_10121) );
NOR2_X2 inst_3348 ( .ZN(net_5577), .A1(net_5436), .A2(net_5435) );
CLKBUF_X2 inst_17993 ( .A(net_9299), .Z(net_17841) );
AOI22_X2 inst_7888 ( .A2(net_4809), .ZN(net_4543), .B2(net_4388), .B1(net_2600), .A1(net_346) );
NAND2_X2 inst_4848 ( .A2(net_8270), .ZN(net_902), .A1(net_663) );
DFFR_X2 inst_7044 ( .QN(net_7520), .D(net_4896), .CK(net_14501), .RN(x6501) );
CLKBUF_X2 inst_15139 ( .A(net_14318), .Z(net_14987) );
CLKBUF_X2 inst_11906 ( .A(net_11753), .Z(net_11754) );
NAND2_X2 inst_4820 ( .A2(net_6381), .A1(net_6380), .ZN(net_1172) );
SDFF_X2 inst_1684 ( .Q(net_8173), .D(net_8173), .SI(net_2639), .SE(net_2538), .CK(net_17125) );
SDFF_X2 inst_1386 ( .SI(net_7301), .Q(net_7118), .D(net_7118), .SE(net_6278), .CK(net_15913) );
XNOR2_X2 inst_217 ( .ZN(net_1412), .B(net_1411), .A(net_700) );
NAND2_X2 inst_4852 ( .A1(net_6148), .ZN(net_896), .A2(net_550) );
NAND2_X2 inst_4616 ( .A2(net_6144), .ZN(net_2609), .A1(net_2608) );
CLKBUF_X2 inst_9816 ( .A(net_9277), .Z(net_9664) );
CLKBUF_X2 inst_15907 ( .A(net_15754), .Z(net_15755) );
SDFFR_X2 inst_2213 ( .Q(net_7465), .D(net_7465), .SE(net_2863), .CK(net_12197), .SI(x13474), .RN(x6501) );
SDFF_X2 inst_672 ( .Q(net_8417), .D(net_8417), .SI(net_3946), .SE(net_3934), .CK(net_10756) );
SDFF_X2 inst_1471 ( .SI(net_7298), .Q(net_7155), .D(net_7155), .SE(net_6279), .CK(net_18195) );
CLKBUF_X2 inst_15393 ( .A(net_15103), .Z(net_15241) );
CLKBUF_X2 inst_17977 ( .A(net_16092), .Z(net_17825) );
CLKBUF_X2 inst_9610 ( .A(net_9457), .Z(net_9458) );
NAND4_X2 inst_3826 ( .A1(net_7210), .ZN(net_2644), .A2(net_2643), .A4(net_2642), .A3(net_1619) );
DFFR_X1 inst_7523 ( .D(net_1295), .Q(net_300), .CK(net_16607), .RN(x6501) );
INV_X2 inst_6471 ( .A(net_7418), .ZN(net_570) );
SDFF_X2 inst_1525 ( .Q(net_7897), .D(net_7897), .SI(net_2749), .SE(net_2543), .CK(net_14415) );
NOR4_X2 inst_3230 ( .ZN(net_2109), .A4(net_1852), .A1(net_505), .A2(x13263), .A3(x13234) );
CLKBUF_X2 inst_11820 ( .A(net_11667), .Z(net_11668) );
CLKBUF_X2 inst_9538 ( .A(net_9385), .Z(net_9386) );
NOR3_X2 inst_3281 ( .ZN(net_2723), .A1(net_2400), .A2(net_2389), .A3(net_2319) );
SDFF_X2 inst_703 ( .Q(net_8422), .D(net_8422), .SI(net_3959), .SE(net_3934), .CK(net_10152) );
CLKBUF_X2 inst_11125 ( .A(net_10972), .Z(net_10973) );
SDFFR_X2 inst_2546 ( .Q(net_6387), .D(net_6387), .SE(net_2147), .SI(net_2127), .CK(net_18243), .RN(x6501) );
CLKBUF_X2 inst_9474 ( .A(net_9318), .Z(net_9322) );
DFFR_X2 inst_7177 ( .QN(net_9013), .D(net_2852), .CK(net_11145), .RN(x6501) );
NAND2_X2 inst_4693 ( .ZN(net_1905), .A2(net_1904), .A1(net_1522) );
CLKBUF_X2 inst_9882 ( .A(net_9729), .Z(net_9730) );
CLKBUF_X2 inst_11112 ( .A(net_10305), .Z(net_10960) );
CLKBUF_X2 inst_12504 ( .A(net_12351), .Z(net_12352) );
CLKBUF_X2 inst_10449 ( .A(net_10296), .Z(net_10297) );
CLKBUF_X2 inst_15737 ( .A(net_15584), .Z(net_15585) );
CLKBUF_X2 inst_14289 ( .A(net_13895), .Z(net_14137) );
CLKBUF_X2 inst_14786 ( .A(net_14633), .Z(net_14634) );
INV_X2 inst_6539 ( .ZN(net_800), .A(net_212) );
SDFF_X2 inst_1067 ( .D(net_7336), .SI(net_6545), .Q(net_6545), .SE(net_3086), .CK(net_9474) );
CLKBUF_X2 inst_12966 ( .A(net_11670), .Z(net_12814) );
DFFR_X1 inst_7411 ( .D(net_5697), .CK(net_16765), .RN(x6501), .Q(x534) );
NAND2_X2 inst_4787 ( .A1(net_2652), .A2(net_1705), .ZN(net_1533) );
CLKBUF_X2 inst_11970 ( .A(net_11817), .Z(net_11818) );
CLKBUF_X2 inst_9735 ( .A(net_9582), .Z(net_9583) );
CLKBUF_X2 inst_9231 ( .A(net_9078), .Z(net_9079) );
SDFF_X2 inst_1824 ( .D(net_7273), .SI(net_6850), .Q(net_6850), .SE(net_6282), .CK(net_14123) );
SDFF_X2 inst_1214 ( .Q(net_7966), .D(net_7966), .SE(net_2755), .SI(net_2717), .CK(net_17037) );
CLKBUF_X2 inst_18580 ( .A(net_14140), .Z(net_18428) );
AOI22_X2 inst_8121 ( .B1(net_8082), .A1(net_7742), .B2(net_6108), .A2(net_6096), .ZN(net_4028) );
CLKBUF_X2 inst_15151 ( .A(net_14998), .Z(net_14999) );
CLKBUF_X2 inst_16197 ( .A(net_11656), .Z(net_16045) );
SDFF_X2 inst_1417 ( .SI(net_7292), .Q(net_7109), .D(net_7109), .SE(net_6278), .CK(net_14925) );
CLKBUF_X2 inst_18510 ( .A(net_15101), .Z(net_18358) );
CLKBUF_X2 inst_11103 ( .A(net_10950), .Z(net_10951) );
CLKBUF_X2 inst_11887 ( .A(net_11439), .Z(net_11735) );
CLKBUF_X2 inst_17803 ( .A(net_17650), .Z(net_17651) );
NOR2_X4 inst_3335 ( .A1(net_6251), .A2(net_6062), .ZN(net_2214) );
OAI21_X2 inst_3073 ( .ZN(net_4223), .A(net_4222), .B2(net_4221), .B1(net_913) );
SDFF_X2 inst_1980 ( .D(net_7293), .SI(net_7030), .Q(net_7030), .SE(net_6277), .CK(net_18351) );
CLKBUF_X2 inst_10488 ( .A(net_10181), .Z(net_10336) );
CLKBUF_X2 inst_17922 ( .A(net_16720), .Z(net_17770) );
CLKBUF_X2 inst_16638 ( .A(net_12124), .Z(net_16486) );
CLKBUF_X2 inst_16792 ( .A(net_15861), .Z(net_16640) );
INV_X4 inst_5868 ( .A(net_8910), .ZN(net_4732) );
OR2_X2 inst_2885 ( .ZN(net_1874), .A2(net_1785), .A1(net_1521) );
CLKBUF_X2 inst_9325 ( .A(net_9172), .Z(net_9173) );
NAND2_X2 inst_4795 ( .ZN(net_3190), .A1(net_1480), .A2(net_1479) );
SDFFR_X2 inst_2632 ( .Q(net_7394), .D(net_7394), .SE(net_1136), .CK(net_15792), .RN(x6501), .SI(x4489) );
SDFFR_X2 inst_2221 ( .Q(net_7449), .D(net_7449), .SE(net_2863), .CK(net_12813), .SI(x13586), .RN(x6501) );
CLKBUF_X2 inst_10446 ( .A(net_9933), .Z(net_10294) );
SDFFS_X2 inst_2082 ( .SI(net_7380), .SE(net_2794), .Q(net_169), .D(net_169), .CK(net_17731), .SN(x6501) );
CLKBUF_X2 inst_12469 ( .A(net_11908), .Z(net_12317) );
CLKBUF_X2 inst_15028 ( .A(net_14325), .Z(net_14876) );
CLKBUF_X2 inst_12907 ( .A(net_12754), .Z(net_12755) );
CLKBUF_X2 inst_15299 ( .A(net_15146), .Z(net_15147) );
CLKBUF_X2 inst_17197 ( .A(net_17044), .Z(net_17045) );
CLKBUF_X2 inst_16204 ( .A(net_13996), .Z(net_16052) );
CLKBUF_X2 inst_13004 ( .A(net_12033), .Z(net_12852) );
SDFF_X2 inst_692 ( .Q(net_8879), .D(net_8879), .SI(net_3941), .SE(net_3936), .CK(net_12879) );
DFF_X1 inst_6800 ( .Q(net_8247), .D(net_4433), .CK(net_13583) );
DFFS_X2 inst_6897 ( .Q(net_6318), .D(net_2638), .CK(net_17455), .SN(x6501) );
CLKBUF_X2 inst_14819 ( .A(net_10186), .Z(net_14667) );
SDFF_X2 inst_1517 ( .Q(net_7884), .D(net_7884), .SI(net_2584), .SE(net_2543), .CK(net_18388) );
CLKBUF_X2 inst_17245 ( .A(net_14611), .Z(net_17093) );
INV_X4 inst_5480 ( .ZN(net_2206), .A(net_737) );
XOR2_X1 inst_70 ( .A(net_3901), .Z(net_3588), .B(net_3587) );
CLKBUF_X2 inst_10529 ( .A(net_10376), .Z(net_10377) );
DFFS_X1 inst_6915 ( .QN(net_6797), .D(net_4723), .CK(net_9551), .SN(x6501) );
CLKBUF_X2 inst_15662 ( .A(net_15509), .Z(net_15510) );
CLKBUF_X2 inst_14161 ( .A(net_14008), .Z(net_14009) );
CLKBUF_X2 inst_15987 ( .A(net_15834), .Z(net_15835) );
INV_X4 inst_6028 ( .ZN(net_505), .A(x13252) );
NAND4_X2 inst_3768 ( .ZN(net_4253), .A1(net_3779), .A2(net_3778), .A3(net_3777), .A4(net_3776) );
CLKBUF_X2 inst_16757 ( .A(net_10508), .Z(net_16605) );
NAND2_X2 inst_4207 ( .ZN(net_5288), .A2(net_5172), .A1(net_5048) );
AND2_X4 inst_9058 ( .A2(net_3325), .ZN(net_3321), .A1(net_3320) );
CLKBUF_X2 inst_11308 ( .A(net_11155), .Z(net_11156) );
INV_X2 inst_6218 ( .ZN(net_5492), .A(net_5357) );
CLKBUF_X2 inst_18550 ( .A(net_11989), .Z(net_18398) );
CLKBUF_X2 inst_13306 ( .A(net_13153), .Z(net_13154) );
OR2_X4 inst_2848 ( .A2(net_4407), .ZN(net_4391), .A1(net_4320) );
CLKBUF_X2 inst_12686 ( .A(net_12533), .Z(net_12534) );
CLKBUF_X2 inst_15181 ( .A(net_15028), .Z(net_15029) );
CLKBUF_X2 inst_18922 ( .A(net_9450), .Z(net_18770) );
CLKBUF_X2 inst_13866 ( .A(net_11602), .Z(net_13714) );
NOR2_X2 inst_3593 ( .ZN(net_2556), .A2(net_833), .A1(x12810) );
CLKBUF_X2 inst_16504 ( .A(net_16351), .Z(net_16352) );
AOI22_X2 inst_8529 ( .B1(net_6723), .A1(net_6690), .B2(net_6202), .A2(net_3520), .ZN(net_3411) );
DFFR_X1 inst_7509 ( .Q(net_6339), .D(net_6338), .CK(net_16951), .RN(x6501) );
OAI211_X4 inst_3176 ( .B(net_6172), .ZN(net_6100), .C1(net_2482), .A(net_2474), .C2(net_1028) );
CLKBUF_X2 inst_15985 ( .A(net_10544), .Z(net_15833) );
CLKBUF_X2 inst_14830 ( .A(net_14677), .Z(net_14678) );
CLKBUF_X2 inst_12655 ( .A(net_12502), .Z(net_12503) );
CLKBUF_X2 inst_13889 ( .A(net_9484), .Z(net_13737) );
CLKBUF_X2 inst_17358 ( .A(net_17205), .Z(net_17206) );
CLKBUF_X2 inst_13730 ( .A(net_12817), .Z(net_13578) );
CLKBUF_X2 inst_10821 ( .A(net_10668), .Z(net_10669) );
SDFF_X2 inst_1150 ( .SI(net_7331), .Q(net_6606), .D(net_6606), .SE(net_3069), .CK(net_11644) );
CLKBUF_X2 inst_17305 ( .A(net_17152), .Z(net_17153) );
MUX2_X2 inst_4914 ( .A(net_6331), .S(net_6330), .Z(net_5933), .B(x4254) );
CLKBUF_X2 inst_18086 ( .A(net_17933), .Z(net_17934) );
CLKBUF_X2 inst_17789 ( .A(net_17636), .Z(net_17637) );
CLKBUF_X2 inst_11020 ( .A(net_10867), .Z(net_10868) );
CLKBUF_X2 inst_11355 ( .A(net_11202), .Z(net_11203) );
CLKBUF_X2 inst_16815 ( .A(net_16662), .Z(net_16663) );
CLKBUF_X2 inst_11770 ( .A(net_9550), .Z(net_11618) );
AOI221_X4 inst_8715 ( .C1(net_7940), .B1(net_7838), .C2(net_6103), .ZN(net_6058), .B2(net_4398), .A(net_4285) );
NAND2_X2 inst_4535 ( .A1(net_3378), .ZN(net_3376), .A2(net_3371) );
CLKBUF_X2 inst_14810 ( .A(net_14657), .Z(net_14658) );
NAND2_X2 inst_4499 ( .A2(net_6272), .ZN(net_4624), .A1(net_1897) );
CLKBUF_X2 inst_12852 ( .A(net_9807), .Z(net_12700) );
DFF_X1 inst_6825 ( .Q(net_8238), .D(net_4442), .CK(net_14451) );
CLKBUF_X2 inst_10979 ( .A(net_10826), .Z(net_10827) );
AOI222_X1 inst_8704 ( .ZN(net_2353), .B1(net_2352), .B2(net_2334), .C2(net_2333), .A2(net_2014), .A1(net_1451), .C1(net_1450) );
CLKBUF_X2 inst_12783 ( .A(net_9698), .Z(net_12631) );
INV_X4 inst_5508 ( .A(net_2935), .ZN(net_858) );
CLKBUF_X2 inst_12661 ( .A(net_12508), .Z(net_12509) );
AOI222_X1 inst_8611 ( .B2(net_6771), .B1(net_5835), .A2(net_5830), .C2(net_5824), .ZN(net_5802), .A1(net_2925), .C1(net_2143) );
SDFF_X2 inst_658 ( .Q(net_8431), .D(net_8431), .SI(net_3942), .SE(net_3934), .CK(net_12610) );
INV_X2 inst_6190 ( .ZN(net_5738), .A(net_5737) );
AOI22_X2 inst_7779 ( .B1(net_6969), .A1(net_6929), .A2(net_5443), .B2(net_5442), .ZN(net_5287) );
CLKBUF_X2 inst_12192 ( .A(net_12039), .Z(net_12040) );
CLKBUF_X2 inst_17728 ( .A(net_16986), .Z(net_17576) );
NAND2_X2 inst_4520 ( .ZN(net_3576), .A2(net_3573), .A1(net_3566) );
DFFR_X2 inst_7227 ( .QN(net_8966), .D(net_2286), .CK(net_13593), .RN(x6501) );
CLKBUF_X2 inst_15090 ( .A(net_11984), .Z(net_14938) );
CLKBUF_X2 inst_9626 ( .A(net_9473), .Z(net_9474) );
CLKBUF_X2 inst_11391 ( .A(net_11238), .Z(net_11239) );
CLKBUF_X2 inst_13581 ( .A(net_12688), .Z(net_13429) );
SDFFR_X2 inst_2128 ( .SI(net_7192), .Q(net_7192), .D(net_6443), .SE(net_4362), .CK(net_13569), .RN(x6501) );
CLKBUF_X2 inst_10452 ( .A(net_10299), .Z(net_10300) );
DFFR_X1 inst_7384 ( .D(net_5847), .CK(net_13907), .RN(x6501), .Q(x608) );
CLKBUF_X2 inst_14472 ( .A(net_10197), .Z(net_14320) );
CLKBUF_X2 inst_10086 ( .A(net_9156), .Z(net_9934) );
CLKBUF_X2 inst_9887 ( .A(net_9734), .Z(net_9735) );
CLKBUF_X2 inst_18066 ( .A(net_17913), .Z(net_17914) );
CLKBUF_X2 inst_11385 ( .A(net_9917), .Z(net_11233) );
AOI22_X2 inst_8289 ( .B1(net_8841), .A1(net_8360), .A2(net_6265), .B2(net_6253), .ZN(net_3753) );
CLKBUF_X2 inst_9313 ( .A(net_9160), .Z(net_9161) );
CLKBUF_X2 inst_10833 ( .A(net_9870), .Z(net_10681) );
NAND2_X2 inst_4455 ( .A2(net_4962), .ZN(net_4960), .A1(net_3252) );
CLKBUF_X2 inst_11402 ( .A(net_11249), .Z(net_11250) );
AOI22_X2 inst_7911 ( .B1(net_8974), .B2(net_5456), .ZN(net_4503), .A2(net_4501), .A1(net_2693) );
CLKBUF_X2 inst_17236 ( .A(net_9387), .Z(net_17084) );
AOI22_X2 inst_7907 ( .A2(net_5538), .ZN(net_4519), .B1(net_4518), .B2(net_4388), .A1(net_421) );
SDFF_X2 inst_929 ( .SI(net_8724), .Q(net_8724), .SE(net_6195), .D(net_3957), .CK(net_12322) );
SDFF_X2 inst_1397 ( .Q(net_8017), .D(net_8017), .SI(net_2658), .SE(net_2545), .CK(net_18064) );
CLKBUF_X2 inst_17327 ( .A(net_17174), .Z(net_17175) );
NOR3_X2 inst_3303 ( .ZN(net_1741), .A1(net_1740), .A3(net_1739), .A2(net_737) );
CLKBUF_X2 inst_13115 ( .A(net_12962), .Z(net_12963) );
INV_X2 inst_6181 ( .ZN(net_5860), .A(net_5815) );
CLKBUF_X2 inst_19166 ( .A(net_19013), .Z(net_19014) );
CLKBUF_X2 inst_12938 ( .A(net_12785), .Z(net_12786) );
INV_X2 inst_6478 ( .ZN(net_887), .A(net_214) );
SDFF_X2 inst_1938 ( .SI(net_8071), .Q(net_8071), .D(net_2639), .SE(net_2508), .CK(net_17113) );
CLKBUF_X2 inst_11870 ( .A(net_11717), .Z(net_11718) );
CLKBUF_X2 inst_9435 ( .A(net_9247), .Z(net_9283) );
DFFS_X2 inst_6888 ( .Q(net_6484), .D(net_2898), .CK(net_9090), .SN(x6501) );
CLKBUF_X2 inst_16020 ( .A(net_15867), .Z(net_15868) );
SDFFS_X2 inst_2095 ( .SI(net_6838), .Q(net_6838), .SE(net_2146), .D(net_1217), .CK(net_18667), .SN(x6501) );
CLKBUF_X2 inst_15659 ( .A(net_15506), .Z(net_15507) );
CLKBUF_X2 inst_18848 ( .A(net_18695), .Z(net_18696) );
CLKBUF_X2 inst_19193 ( .A(net_19040), .Z(net_19041) );
INV_X4 inst_5794 ( .A(net_6294), .ZN(net_1198) );
CLKBUF_X2 inst_14103 ( .A(net_13950), .Z(net_13951) );
AOI21_X2 inst_8896 ( .B2(net_5871), .ZN(net_5789), .A(net_5788), .B1(net_2640) );
INV_X4 inst_5652 ( .A(net_7397), .ZN(net_943) );
AOI22_X2 inst_8262 ( .B1(net_8874), .A1(net_8319), .B2(net_6252), .A2(net_4345), .ZN(net_3776) );
INV_X4 inst_5631 ( .A(net_8940), .ZN(net_2620) );
SDFF_X2 inst_683 ( .Q(net_8685), .D(net_8685), .SI(net_3958), .SE(net_3935), .CK(net_10998) );
CLKBUF_X2 inst_11813 ( .A(net_11660), .Z(net_11661) );
CLKBUF_X2 inst_17144 ( .A(net_16991), .Z(net_16992) );
AND2_X4 inst_9094 ( .A1(net_2501), .ZN(net_2483), .A2(net_2197) );
CLKBUF_X2 inst_9411 ( .A(net_9258), .Z(net_9259) );
AOI221_X4 inst_8720 ( .B1(net_8720), .C1(net_8498), .B2(net_4350), .C2(net_4349), .ZN(net_4347), .A(net_4260) );
CLKBUF_X2 inst_17418 ( .A(net_17265), .Z(net_17266) );
CLKBUF_X2 inst_12103 ( .A(net_11950), .Z(net_11951) );
INV_X4 inst_5893 ( .A(net_6298), .ZN(net_2690) );
NAND3_X4 inst_3881 ( .A2(net_5980), .A1(net_1561), .ZN(net_1530), .A3(net_1529) );
CLKBUF_X2 inst_18730 ( .A(net_18577), .Z(net_18578) );
NAND2_X2 inst_4778 ( .ZN(net_1785), .A1(net_1703), .A2(net_1614) );
CLKBUF_X2 inst_14580 ( .A(net_14427), .Z(net_14428) );
CLKBUF_X2 inst_17884 ( .A(net_17030), .Z(net_17732) );
INV_X4 inst_5325 ( .ZN(net_1618), .A(net_1520) );
NAND2_X2 inst_4576 ( .A1(net_7172), .A2(net_3035), .ZN(net_3026) );
SDFF_X2 inst_747 ( .Q(net_8790), .D(net_8790), .SI(net_3945), .SE(net_3879), .CK(net_13333) );
CLKBUF_X2 inst_15493 ( .A(net_13188), .Z(net_15341) );
HA_X1 inst_6685 ( .S(net_3011), .CO(net_3010), .A(net_3009), .B(net_2865) );
AND2_X4 inst_9070 ( .ZN(net_6138), .A1(net_3250), .A2(net_3215) );
NAND4_X2 inst_3806 ( .ZN(net_3620), .A1(net_3463), .A2(net_3462), .A3(net_3461), .A4(net_3460) );
CLKBUF_X2 inst_18594 ( .A(net_18441), .Z(net_18442) );
NAND2_X2 inst_4486 ( .A2(net_5267), .ZN(net_4492), .A1(net_174) );
CLKBUF_X2 inst_15964 ( .A(net_13708), .Z(net_15812) );
CLKBUF_X2 inst_12893 ( .A(net_12740), .Z(net_12741) );
CLKBUF_X2 inst_17747 ( .A(net_17594), .Z(net_17595) );
CLKBUF_X2 inst_11362 ( .A(net_11209), .Z(net_11210) );
CLKBUF_X2 inst_14946 ( .A(net_14793), .Z(net_14794) );
SDFFR_X1 inst_2775 ( .D(net_7385), .Q(net_7282), .SI(net_1955), .SE(net_1327), .CK(net_15375), .RN(x6501) );
INV_X4 inst_5589 ( .A(net_7381), .ZN(net_654) );
CLKBUF_X2 inst_15324 ( .A(net_15171), .Z(net_15172) );
CLKBUF_X2 inst_19040 ( .A(net_18887), .Z(net_18888) );
CLKBUF_X2 inst_12334 ( .A(net_12181), .Z(net_12182) );
XNOR2_X2 inst_305 ( .B(net_1864), .ZN(net_968), .A(net_504) );
DFF_X1 inst_6795 ( .QN(net_8242), .D(net_4438), .CK(net_17597) );
CLKBUF_X2 inst_13516 ( .A(net_13363), .Z(net_13364) );
SDFF_X2 inst_1595 ( .Q(net_8128), .D(net_8128), .SI(net_2575), .SE(net_2541), .CK(net_15993) );
AOI22_X2 inst_7881 ( .B1(net_7195), .A2(net_6446), .B2(net_5655), .A1(net_5654), .ZN(net_4550) );
INV_X4 inst_5651 ( .A(net_6470), .ZN(net_980) );
AOI22_X2 inst_7867 ( .B2(net_5609), .A2(net_5267), .ZN(net_4574), .B1(net_381), .A1(net_185) );
CLKBUF_X2 inst_15922 ( .A(net_15769), .Z(net_15770) );
CLKBUF_X2 inst_10926 ( .A(net_10773), .Z(net_10774) );
CLKBUF_X2 inst_13578 ( .A(net_13425), .Z(net_13426) );
CLKBUF_X2 inst_12319 ( .A(net_12166), .Z(net_12167) );
AOI22_X2 inst_8079 ( .B1(net_7910), .A1(net_7808), .B2(net_6103), .A2(net_4398), .ZN(net_4066) );
INV_X2 inst_6585 ( .A(net_7507), .ZN(net_477) );
CLKBUF_X2 inst_13069 ( .A(net_12916), .Z(net_12917) );
CLKBUF_X2 inst_15595 ( .A(net_11985), .Z(net_15443) );
AOI22_X2 inst_7774 ( .B1(net_6964), .A1(net_6924), .A2(net_5443), .B2(net_5442), .ZN(net_5307) );
SDFF_X2 inst_963 ( .SI(net_7321), .Q(net_6728), .D(net_6728), .SE(net_3124), .CK(net_12126) );
CLKBUF_X2 inst_17986 ( .A(net_17163), .Z(net_17834) );
CLKBUF_X2 inst_16787 ( .A(net_16634), .Z(net_16635) );
SDFF_X2 inst_1614 ( .Q(net_8146), .D(net_8146), .SI(net_2721), .SE(net_2538), .CK(net_15762) );
SDFF_X2 inst_1502 ( .SI(net_7860), .Q(net_7860), .D(net_2718), .SE(net_2558), .CK(net_14917) );
INV_X4 inst_5436 ( .A(net_7212), .ZN(net_825) );
INV_X4 inst_6115 ( .ZN(net_1916), .A(net_262) );
NAND2_X2 inst_4091 ( .ZN(net_5447), .A1(net_5251), .A2(net_5018) );
CLKBUF_X2 inst_16732 ( .A(net_16579), .Z(net_16580) );
DFFR_X2 inst_6989 ( .D(net_5896), .CK(net_11490), .RN(x6501), .Q(x2693) );
DFF_X1 inst_6807 ( .Q(net_8224), .D(net_4421), .CK(net_16554) );
CLKBUF_X2 inst_15854 ( .A(net_15701), .Z(net_15702) );
SDFF_X2 inst_1568 ( .Q(net_8112), .D(net_8112), .SI(net_2721), .SE(net_2541), .CK(net_15829) );
CLKBUF_X2 inst_11439 ( .A(net_11286), .Z(net_11287) );
INV_X2 inst_6177 ( .ZN(net_5911), .A(net_5866) );
AOI22_X2 inst_8487 ( .B1(net_6611), .A1(net_6578), .A2(net_6257), .B2(net_6110), .ZN(net_3453) );
NOR2_X2 inst_3366 ( .ZN(net_5559), .A1(net_5364), .A2(net_5363) );
SDFF_X2 inst_873 ( .Q(net_8584), .D(net_8584), .SI(net_3953), .SE(net_3878), .CK(net_10225) );
CLKBUF_X2 inst_9258 ( .A(net_9105), .Z(net_9106) );
CLKBUF_X2 inst_12223 ( .A(net_10357), .Z(net_12071) );
INV_X2 inst_6454 ( .A(net_6364), .ZN(net_2143) );
CLKBUF_X2 inst_13439 ( .A(net_10784), .Z(net_13287) );
CLKBUF_X2 inst_10022 ( .A(net_9869), .Z(net_9870) );
CLKBUF_X2 inst_10164 ( .A(net_10011), .Z(net_10012) );
CLKBUF_X2 inst_16614 ( .A(net_16461), .Z(net_16462) );
AOI22_X2 inst_8563 ( .A1(net_2694), .A2(net_2334), .B2(net_2333), .ZN(net_2330), .B1(net_1846) );
NAND4_X2 inst_3767 ( .A3(net_6065), .A1(net_6064), .ZN(net_4254), .A2(net_3784), .A4(net_3783) );
CLKBUF_X2 inst_10282 ( .A(net_10129), .Z(net_10130) );
AOI221_X2 inst_8839 ( .C1(net_8183), .B1(net_7673), .C2(net_6099), .ZN(net_5991), .B2(net_4399), .A(net_4283) );
NAND2_X2 inst_4431 ( .A1(net_6869), .A2(net_5016), .ZN(net_4996) );
AOI222_X1 inst_8679 ( .B1(net_6752), .A1(net_6460), .ZN(net_3297), .A2(net_3296), .B2(net_3295), .C2(net_3294), .C1(net_2949) );
NOR2_X2 inst_3371 ( .ZN(net_5554), .A1(net_5344), .A2(net_5343) );
OAI21_X2 inst_3052 ( .B2(net_8233), .B1(net_4850), .ZN(net_4759), .A(net_2593) );
CLKBUF_X2 inst_15920 ( .A(net_15767), .Z(net_15768) );
DFFR_X2 inst_6982 ( .QN(net_5966), .D(net_5905), .CK(net_9342), .RN(x6501) );
CLKBUF_X2 inst_17210 ( .A(net_17057), .Z(net_17058) );
CLKBUF_X2 inst_16942 ( .A(net_16789), .Z(net_16790) );
OAI22_X4 inst_2907 ( .ZN(net_6134), .B2(net_4512), .A1(net_4472), .A2(net_4407), .B1(net_4391) );
CLKBUF_X2 inst_13548 ( .A(net_13395), .Z(net_13396) );
NAND2_X2 inst_4072 ( .A2(net_6789), .A1(net_5775), .ZN(net_5774) );
INV_X4 inst_5901 ( .A(net_7349), .ZN(net_638) );
OAI21_X2 inst_3000 ( .B2(net_5902), .ZN(net_5893), .A(net_5817), .B1(net_618) );
SDFF_X2 inst_1163 ( .SI(net_7317), .Q(net_6592), .D(net_6592), .SE(net_3069), .CK(net_11993) );
CLKBUF_X2 inst_9668 ( .A(net_9373), .Z(net_9516) );
CLKBUF_X2 inst_10641 ( .A(net_10036), .Z(net_10489) );
AOI22_X2 inst_8282 ( .B1(net_8692), .A1(net_8655), .B2(net_6109), .A2(net_3857), .ZN(net_3759) );
CLKBUF_X2 inst_18399 ( .A(net_10980), .Z(net_18247) );
NOR4_X2 inst_3239 ( .ZN(net_1718), .A2(net_1362), .A3(net_1250), .A1(net_793), .A4(net_784) );
SDFFR_X2 inst_2314 ( .SE(net_2260), .Q(net_370), .D(net_370), .CK(net_9174), .RN(x6501), .SI(x1667) );
CLKBUF_X2 inst_12885 ( .A(net_10180), .Z(net_12733) );
OR3_X2 inst_2812 ( .A3(net_5957), .ZN(net_1525), .A1(net_1524), .A2(net_1523) );
NAND2_X2 inst_4743 ( .ZN(net_2712), .A2(net_1586), .A1(net_922) );
CLKBUF_X2 inst_15607 ( .A(net_9810), .Z(net_15455) );
OAI211_X2 inst_3197 ( .ZN(net_3035), .C2(net_2892), .A(net_2399), .B(net_2086), .C1(net_1368) );
NAND2_X2 inst_4651 ( .A1(net_6115), .ZN(net_5044), .A2(net_2580) );
CLKBUF_X2 inst_10126 ( .A(net_9973), .Z(net_9974) );
CLKBUF_X2 inst_13640 ( .A(net_13487), .Z(net_13488) );
AOI22_X2 inst_8006 ( .B1(net_8011), .A1(net_7977), .B2(net_6102), .A2(net_6097), .ZN(net_4128) );
CLKBUF_X2 inst_14988 ( .A(net_14835), .Z(net_14836) );
SDFF_X2 inst_1083 ( .D(net_7336), .SI(net_6512), .Q(net_6512), .SE(net_3071), .CK(net_11680) );
NAND2_X2 inst_4073 ( .A2(net_6790), .A1(net_5775), .ZN(net_5773) );
INV_X4 inst_6123 ( .A(net_5979), .ZN(x3712) );
SDFFR_X2 inst_2466 ( .SE(net_2683), .D(net_2571), .SI(net_438), .Q(net_438), .CK(net_14542), .RN(x6501) );
CLKBUF_X2 inst_11979 ( .A(net_11826), .Z(net_11827) );
CLKBUF_X2 inst_11877 ( .A(net_9710), .Z(net_11725) );
CLKBUF_X2 inst_12070 ( .A(net_11917), .Z(net_11918) );
CLKBUF_X2 inst_13615 ( .A(net_13462), .Z(net_13463) );
SDFF_X2 inst_696 ( .Q(net_8444), .D(net_8444), .SI(net_3948), .SE(net_3934), .CK(net_13407) );
CLKBUF_X2 inst_9719 ( .A(net_9146), .Z(net_9567) );
CLKBUF_X2 inst_11890 ( .A(net_11737), .Z(net_11738) );
CLKBUF_X2 inst_15555 ( .A(net_15402), .Z(net_15403) );
CLKBUF_X2 inst_10755 ( .A(net_10602), .Z(net_10603) );
CLKBUF_X2 inst_12059 ( .A(net_10068), .Z(net_11907) );
INV_X8 inst_5055 ( .ZN(net_6274), .A(net_6261) );
INV_X4 inst_6128 ( .A(net_6359), .ZN(net_481) );
CLKBUF_X2 inst_10778 ( .A(net_9401), .Z(net_10626) );
NAND3_X2 inst_3969 ( .ZN(net_2548), .A2(net_2279), .A1(net_2278), .A3(net_2181) );
CLKBUF_X2 inst_11712 ( .A(net_10159), .Z(net_11560) );
SDFFR_X2 inst_2363 ( .SI(net_7366), .SE(net_2732), .D(net_1817), .QN(net_270), .CK(net_16120), .RN(x6501) );
CLKBUF_X2 inst_9909 ( .A(net_9756), .Z(net_9757) );
INV_X4 inst_6014 ( .A(net_5966), .ZN(x3122) );
INV_X2 inst_6257 ( .ZN(net_4695), .A(net_4665) );
NAND2_X4 inst_4029 ( .A2(net_6218), .A1(net_6183), .ZN(net_5989) );
SDFF_X2 inst_1629 ( .Q(net_8174), .D(net_8174), .SI(net_2715), .SE(net_2538), .CK(net_14266) );
CLKBUF_X2 inst_16999 ( .A(net_13865), .Z(net_16847) );
CLKBUF_X2 inst_17061 ( .A(net_16908), .Z(net_16909) );
CLKBUF_X2 inst_15583 ( .A(net_15430), .Z(net_15431) );
NOR2_X2 inst_3424 ( .ZN(net_3094), .A2(net_3093), .A1(net_2983) );
CLKBUF_X2 inst_17840 ( .A(net_17687), .Z(net_17688) );
CLKBUF_X2 inst_12138 ( .A(net_9126), .Z(net_11986) );
CLKBUF_X2 inst_13923 ( .A(net_12620), .Z(net_13771) );
CLKBUF_X2 inst_15895 ( .A(net_15742), .Z(net_15743) );
SDFFR_X2 inst_2580 ( .D(net_7378), .QN(net_7238), .SI(net_1956), .SE(net_1379), .CK(net_17518), .RN(x6501) );
CLKBUF_X2 inst_11342 ( .A(net_11189), .Z(net_11190) );
CLKBUF_X2 inst_16799 ( .A(net_16646), .Z(net_16647) );
CLKBUF_X2 inst_14213 ( .A(net_11651), .Z(net_14061) );
CLKBUF_X2 inst_12268 ( .A(net_12115), .Z(net_12116) );
CLKBUF_X2 inst_17103 ( .A(net_14583), .Z(net_16951) );
INV_X4 inst_5840 ( .A(net_8258), .ZN(net_3029) );
CLKBUF_X2 inst_15290 ( .A(net_15137), .Z(net_15138) );
SDFF_X2 inst_2054 ( .SI(net_7802), .Q(net_7802), .D(net_2704), .SE(net_2459), .CK(net_16961) );
CLKBUF_X2 inst_12216 ( .A(net_12063), .Z(net_12064) );
CLKBUF_X2 inst_13448 ( .A(net_11207), .Z(net_13296) );
SDFF_X2 inst_1259 ( .Q(net_8100), .D(net_8100), .SI(net_2712), .SE(net_2707), .CK(net_13797) );
CLKBUF_X2 inst_18216 ( .A(net_18063), .Z(net_18064) );
CLKBUF_X2 inst_16148 ( .A(net_15995), .Z(net_15996) );
AOI22_X2 inst_7821 ( .B1(net_7511), .A2(net_5535), .B2(net_5260), .ZN(net_4703), .A1(net_470) );
SDFF_X2 inst_1796 ( .D(net_7293), .SI(net_6870), .Q(net_6870), .SE(net_6282), .CK(net_17684) );
CLKBUF_X2 inst_10702 ( .A(net_10549), .Z(net_10550) );
CLKBUF_X2 inst_18573 ( .A(net_12892), .Z(net_18421) );
CLKBUF_X2 inst_12318 ( .A(net_12165), .Z(net_12166) );
SDFF_X2 inst_535 ( .Q(net_8857), .D(net_8857), .SI(net_3965), .SE(net_3936), .CK(net_11093) );
CLKBUF_X2 inst_11341 ( .A(net_11188), .Z(net_11189) );
CLKBUF_X2 inst_12970 ( .A(net_12817), .Z(net_12818) );
AOI22_X2 inst_7853 ( .A2(net_5595), .B2(net_4881), .ZN(net_4654), .A1(net_324), .B1(net_242) );
CLKBUF_X2 inst_10059 ( .A(net_9658), .Z(net_9907) );
CLKBUF_X2 inst_16589 ( .A(net_16436), .Z(net_16437) );
SDFFR_X2 inst_2427 ( .D(net_2674), .SE(net_2313), .SI(net_450), .Q(net_450), .CK(net_16535), .RN(x6501) );
CLKBUF_X2 inst_11670 ( .A(net_11517), .Z(net_11518) );
AOI222_X1 inst_8603 ( .B2(net_6768), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5821), .A1(net_2885), .C1(x3122) );
CLKBUF_X2 inst_10496 ( .A(net_9358), .Z(net_10344) );
NOR3_X2 inst_3317 ( .A2(net_7258), .A3(net_7225), .ZN(net_2084), .A1(net_1802) );
CLKBUF_X2 inst_14616 ( .A(net_12874), .Z(net_14464) );
CLKBUF_X2 inst_17399 ( .A(net_17246), .Z(net_17247) );
INV_X4 inst_6079 ( .A(net_6310), .ZN(net_2729) );
CLKBUF_X2 inst_13245 ( .A(net_13092), .Z(net_13093) );
CLKBUF_X2 inst_11348 ( .A(net_11195), .Z(net_11196) );
DFFR_X2 inst_7206 ( .D(net_2367), .QN(net_219), .CK(net_14725), .RN(x6501) );
OAI21_X2 inst_3168 ( .ZN(net_1528), .B1(net_1527), .B2(net_1526), .A(net_1336) );
NAND4_X2 inst_3855 ( .A1(net_6383), .A3(net_6382), .A4(net_6380), .ZN(net_1260), .A2(net_1258) );
AOI222_X2 inst_8589 ( .B2(net_8247), .B1(net_4891), .C2(net_4889), .ZN(net_4839), .A1(net_4803), .A2(net_3547), .C1(net_3546) );
NOR3_X2 inst_3318 ( .ZN(net_1663), .A1(net_1283), .A3(net_1085), .A2(net_687) );
CLKBUF_X2 inst_10594 ( .A(net_10441), .Z(net_10442) );
CLKBUF_X2 inst_12771 ( .A(net_9797), .Z(net_12619) );
CLKBUF_X2 inst_10299 ( .A(net_9747), .Z(net_10147) );
INV_X4 inst_5176 ( .ZN(net_3948), .A(net_2907) );
CLKBUF_X2 inst_12672 ( .A(net_12519), .Z(net_12520) );
CLKBUF_X2 inst_19145 ( .A(net_18992), .Z(net_18993) );
SDFF_X2 inst_1322 ( .Q(net_7945), .D(net_7945), .SE(net_2755), .SI(net_2655), .CK(net_18568) );
CLKBUF_X2 inst_11862 ( .A(net_11709), .Z(net_11710) );
CLKBUF_X2 inst_16483 ( .A(net_16330), .Z(net_16331) );
CLKBUF_X2 inst_17380 ( .A(net_17227), .Z(net_17228) );
CLKBUF_X2 inst_10954 ( .A(net_9500), .Z(net_10802) );
CLKBUF_X2 inst_14891 ( .A(net_12840), .Z(net_14739) );
CLKBUF_X2 inst_14004 ( .A(net_13851), .Z(net_13852) );
CLKBUF_X2 inst_10712 ( .A(net_10444), .Z(net_10560) );
CLKBUF_X2 inst_14237 ( .A(net_10153), .Z(net_14085) );
CLKBUF_X2 inst_10248 ( .A(net_9932), .Z(net_10096) );
CLKBUF_X2 inst_15471 ( .A(net_15318), .Z(net_15319) );
CLKBUF_X2 inst_17029 ( .A(net_16876), .Z(net_16877) );
AOI22_X2 inst_8379 ( .B1(net_8560), .A1(net_8449), .A2(net_6263), .B2(net_6262), .ZN(net_3669) );
CLKBUF_X2 inst_10156 ( .A(net_10003), .Z(net_10004) );
NOR2_X2 inst_3493 ( .A1(net_3023), .ZN(net_2035), .A2(net_1851) );
CLKBUF_X2 inst_9776 ( .A(net_9623), .Z(net_9624) );
CLKBUF_X2 inst_10413 ( .A(net_9841), .Z(net_10261) );
CLKBUF_X2 inst_13151 ( .A(net_12998), .Z(net_12999) );
NAND2_X2 inst_4622 ( .A2(net_6144), .ZN(net_2597), .A1(net_2596) );
NOR2_X2 inst_3487 ( .A2(net_2400), .ZN(net_2278), .A1(net_2180) );
NOR2_X2 inst_3597 ( .ZN(net_1333), .A1(net_1271), .A2(net_909) );
CLKBUF_X2 inst_11783 ( .A(net_11630), .Z(net_11631) );
CLKBUF_X2 inst_14421 ( .A(net_10216), .Z(net_14269) );
CLKBUF_X2 inst_14555 ( .A(net_14402), .Z(net_14403) );
AOI22_X2 inst_8210 ( .B1(net_8757), .A1(net_8387), .A2(net_3867), .B2(net_3866), .ZN(net_3826) );
CLKBUF_X2 inst_10661 ( .A(net_10508), .Z(net_10509) );
CLKBUF_X2 inst_11757 ( .A(net_11604), .Z(net_11605) );
CLKBUF_X2 inst_13422 ( .A(net_13269), .Z(net_13270) );
SDFFR_X2 inst_2607 ( .D(net_7375), .Q(net_7272), .SI(net_1807), .SE(net_1327), .CK(net_17507), .RN(x6501) );
CLKBUF_X2 inst_16287 ( .A(net_16134), .Z(net_16135) );
AOI22_X2 inst_8133 ( .B1(net_8152), .A1(net_7710), .B2(net_6101), .A2(net_6095), .ZN(net_6030) );
CLKBUF_X2 inst_13893 ( .A(net_13740), .Z(net_13741) );
CLKBUF_X2 inst_11395 ( .A(net_11242), .Z(net_11243) );
AOI22_X2 inst_7791 ( .B2(net_6187), .A2(net_6134), .ZN(net_4807), .A1(net_1399), .B1(net_202) );
SDFFR_X1 inst_2690 ( .SI(net_7554), .SE(net_5043), .CK(net_12746), .RN(x6501), .Q(x3861), .D(x3861) );
AOI222_X1 inst_8689 ( .C2(net_5832), .A2(net_5830), .B2(net_5824), .ZN(net_3280), .A1(net_3102), .B1(net_2135), .C1(x2594) );
CLKBUF_X2 inst_10467 ( .A(net_9649), .Z(net_10315) );
CLKBUF_X2 inst_16167 ( .A(net_9143), .Z(net_16015) );
SDFF_X2 inst_1544 ( .Q(net_7999), .D(net_7999), .SI(net_2749), .SE(net_2542), .CK(net_14411) );
INV_X2 inst_6261 ( .A(net_8240), .ZN(net_4636) );
CLKBUF_X2 inst_9771 ( .A(net_9618), .Z(net_9619) );
OAI21_X2 inst_3148 ( .B2(net_2048), .ZN(net_1989), .A(net_1988), .B1(net_764) );
CLKBUF_X2 inst_17721 ( .A(net_9625), .Z(net_17569) );
NAND2_X2 inst_4761 ( .ZN(net_2293), .A1(net_399), .A2(net_396) );
INV_X4 inst_5180 ( .A(net_3033), .ZN(net_2999) );
OAI21_X2 inst_3026 ( .ZN(net_4958), .A(net_4957), .B2(net_4956), .B1(net_4924) );
DFFS_X1 inst_6952 ( .QN(net_6472), .D(net_3342), .CK(net_15087), .SN(x6501) );
AOI22_X2 inst_8573 ( .A1(net_2546), .B2(net_1919), .A2(net_1918), .ZN(net_1917), .B1(net_1916) );
CLKBUF_X2 inst_17017 ( .A(net_9394), .Z(net_16865) );
NAND4_X2 inst_3639 ( .ZN(net_5025), .A4(net_4769), .A1(net_4698), .A3(net_4696), .A2(net_4667) );
CLKBUF_X2 inst_13646 ( .A(net_13493), .Z(net_13494) );
DFFR_X2 inst_7226 ( .QN(net_9006), .D(net_2236), .CK(net_16290), .RN(x6501) );
AND2_X2 inst_9194 ( .ZN(net_1759), .A1(net_1581), .A2(net_1580) );
CLKBUF_X2 inst_10411 ( .A(net_10258), .Z(net_10259) );
CLKBUF_X2 inst_13130 ( .A(net_12977), .Z(net_12978) );
CLKBUF_X2 inst_14241 ( .A(net_9502), .Z(net_14089) );
CLKBUF_X2 inst_12769 ( .A(net_12616), .Z(net_12617) );
SDFF_X2 inst_752 ( .Q(net_8792), .D(net_8792), .SI(net_3959), .SE(net_3879), .CK(net_13177) );
NOR4_X2 inst_3245 ( .ZN(net_1558), .A4(net_1017), .A3(net_1005), .A1(net_996), .A2(net_954) );
OAI211_X2 inst_3202 ( .C2(net_2652), .ZN(net_2425), .A(net_2424), .B(net_2423), .C1(net_2179) );
NAND2_X2 inst_4279 ( .A1(net_6884), .A2(net_5247), .ZN(net_5181) );
CLKBUF_X2 inst_18125 ( .A(net_9104), .Z(net_17973) );
SDFF_X2 inst_1384 ( .SI(net_7264), .Q(net_7121), .D(net_7121), .SE(net_6279), .CK(net_14372) );
CLKBUF_X2 inst_16116 ( .A(net_15687), .Z(net_15964) );
SDFFR_X2 inst_2118 ( .SI(net_7176), .Q(net_7176), .D(net_6427), .SE(net_4362), .CK(net_13577), .RN(x6501) );
CLKBUF_X2 inst_16112 ( .A(net_15959), .Z(net_15960) );
AOI22_X2 inst_7749 ( .B1(net_6978), .A1(net_6938), .A2(net_5443), .B2(net_5442), .ZN(net_5410) );
CLKBUF_X2 inst_18347 ( .A(net_18194), .Z(net_18195) );
AOI221_X2 inst_8817 ( .C2(net_5535), .B2(net_5260), .A(net_4898), .ZN(net_4710), .B1(net_3236), .C1(net_463) );
INV_X8 inst_5048 ( .A(net_6169), .ZN(net_6168) );
CLKBUF_X2 inst_18866 ( .A(net_18713), .Z(net_18714) );
CLKBUF_X2 inst_11470 ( .A(net_11317), .Z(net_11318) );
CLKBUF_X2 inst_12693 ( .A(net_11228), .Z(net_12541) );
NAND2_X2 inst_4356 ( .A1(net_7122), .A2(net_5166), .ZN(net_5101) );
CLKBUF_X2 inst_18753 ( .A(net_15845), .Z(net_18601) );
CLKBUF_X2 inst_18226 ( .A(net_18073), .Z(net_18074) );
CLKBUF_X2 inst_16761 ( .A(net_16608), .Z(net_16609) );
CLKBUF_X2 inst_11707 ( .A(net_11554), .Z(net_11555) );
CLKBUF_X2 inst_9975 ( .A(net_9822), .Z(net_9823) );
CLKBUF_X2 inst_12250 ( .A(net_9448), .Z(net_12098) );
INV_X4 inst_5329 ( .ZN(net_1607), .A(net_1350) );
SDFFR_X2 inst_2539 ( .QN(net_6375), .SE(net_2147), .SI(net_1960), .D(net_617), .CK(net_18326), .RN(x6501) );
CLKBUF_X2 inst_10141 ( .A(net_9988), .Z(net_9989) );
CLKBUF_X2 inst_13496 ( .A(net_13343), .Z(net_13344) );
OR3_X4 inst_2797 ( .ZN(net_3337), .A3(net_3278), .A1(net_3243), .A2(net_1074) );
NOR2_X2 inst_3431 ( .A2(net_3093), .ZN(net_3078), .A1(net_1187) );
CLKBUF_X2 inst_13193 ( .A(net_12517), .Z(net_13041) );
SDFFS_X2 inst_2085 ( .SI(net_7383), .SE(net_2795), .Q(net_172), .D(net_172), .CK(net_17430), .SN(x6501) );
CLKBUF_X2 inst_17062 ( .A(net_13923), .Z(net_16910) );
CLKBUF_X2 inst_11097 ( .A(net_10944), .Z(net_10945) );
INV_X4 inst_5264 ( .ZN(net_2672), .A(net_1586) );
CLKBUF_X2 inst_12910 ( .A(net_10823), .Z(net_12758) );
DFFR_X2 inst_7069 ( .QN(net_7417), .D(net_4202), .CK(net_12303), .RN(x6501) );
INV_X4 inst_6150 ( .A(net_6164), .ZN(net_6162) );
CLKBUF_X2 inst_14230 ( .A(net_14066), .Z(net_14078) );
SDFF_X2 inst_556 ( .Q(net_8670), .D(net_8670), .SI(net_3977), .SE(net_3935), .CK(net_11091) );
CLKBUF_X2 inst_11779 ( .A(net_11626), .Z(net_11627) );
NAND4_X2 inst_3632 ( .ZN(net_5528), .A2(net_5038), .A4(net_4871), .A3(net_4812), .A1(net_4463) );
INV_X4 inst_5147 ( .A(net_3243), .ZN(net_3242) );
CLKBUF_X2 inst_13758 ( .A(net_13605), .Z(net_13606) );
CLKBUF_X2 inst_12573 ( .A(net_12420), .Z(net_12421) );
CLKBUF_X2 inst_9650 ( .A(net_9497), .Z(net_9498) );
CLKBUF_X2 inst_15641 ( .A(net_15488), .Z(net_15489) );
NOR3_X2 inst_3300 ( .ZN(net_1831), .A3(net_1557), .A1(net_1213), .A2(net_969) );
CLKBUF_X2 inst_16457 ( .A(net_14424), .Z(net_16305) );
CLKBUF_X2 inst_12728 ( .A(net_12575), .Z(net_12576) );
NAND4_X2 inst_3822 ( .ZN(net_3604), .A1(net_3399), .A2(net_3398), .A3(net_3397), .A4(net_3396) );
AOI221_X2 inst_8757 ( .C2(net_5609), .ZN(net_5521), .B2(net_5520), .A(net_5025), .C1(net_356), .B1(net_286) );
CLKBUF_X2 inst_9603 ( .A(net_9059), .Z(net_9451) );
DFFR_X1 inst_7522 ( .D(net_824), .Q(net_298), .CK(net_15216), .RN(x6501) );
NAND2_X2 inst_4593 ( .ZN(net_3928), .A2(net_2845), .A1(net_2799) );
INV_X4 inst_6070 ( .A(net_7492), .ZN(net_4884) );
CLKBUF_X2 inst_17769 ( .A(net_17616), .Z(net_17617) );
NOR3_X2 inst_3307 ( .A3(net_2666), .ZN(net_2204), .A1(net_1338), .A2(net_642) );
SDFF_X2 inst_1587 ( .Q(net_8043), .D(net_8043), .SI(net_2703), .SE(net_2545), .CK(net_14009) );
INV_X4 inst_5452 ( .ZN(net_2397), .A(net_801) );
SDFF_X2 inst_1185 ( .D(net_7339), .SI(net_6581), .Q(net_6581), .SE(net_3070), .CK(net_9601) );
CLKBUF_X2 inst_16262 ( .A(net_16109), .Z(net_16110) );
AOI221_X2 inst_8742 ( .C1(net_8998), .ZN(net_5662), .A(net_5583), .B2(net_5538), .C2(net_5456), .B1(net_427) );
SDFF_X2 inst_457 ( .SI(net_8460), .Q(net_8460), .SE(net_3983), .D(net_3973), .CK(net_12355) );
CLKBUF_X2 inst_13715 ( .A(net_13562), .Z(net_13563) );
CLKBUF_X2 inst_16213 ( .A(net_16060), .Z(net_16061) );
SDFF_X2 inst_1738 ( .Q(net_8207), .D(net_8207), .SI(net_2639), .SE(net_2561), .CK(net_17121) );
OR3_X4 inst_2802 ( .A3(net_6112), .ZN(net_2424), .A1(net_1322), .A2(net_820) );
NAND2_X2 inst_4171 ( .ZN(net_5339), .A2(net_5196), .A1(net_5084) );
CLKBUF_X2 inst_15169 ( .A(net_15016), .Z(net_15017) );
CLKBUF_X2 inst_11276 ( .A(net_11123), .Z(net_11124) );
CLKBUF_X2 inst_16385 ( .A(net_16232), .Z(net_16233) );
DFFR_X2 inst_7204 ( .QN(net_6394), .D(net_2301), .CK(net_15675), .RN(x6501) );
INV_X4 inst_5529 ( .ZN(net_877), .A(net_661) );
CLKBUF_X2 inst_14984 ( .A(net_14831), .Z(net_14832) );
AOI21_X2 inst_8953 ( .A(net_5746), .ZN(net_5659), .B1(net_5474), .B2(net_5457) );
CLKBUF_X2 inst_10250 ( .A(net_10097), .Z(net_10098) );
CLKBUF_X2 inst_16259 ( .A(net_16106), .Z(net_16107) );
INV_X4 inst_6103 ( .A(net_7345), .ZN(net_3258) );
CLKBUF_X2 inst_16953 ( .A(net_16800), .Z(net_16801) );
XNOR2_X2 inst_146 ( .ZN(net_2227), .B(net_2139), .A(net_2138) );
CLKBUF_X2 inst_15588 ( .A(net_13852), .Z(net_15436) );
NAND3_X2 inst_3999 ( .A3(net_7402), .ZN(net_4407), .A1(net_1105), .A2(net_499) );
CLKBUF_X2 inst_18710 ( .A(net_10415), .Z(net_18558) );
CLKBUF_X2 inst_18703 ( .A(net_15760), .Z(net_18551) );
CLKBUF_X2 inst_12501 ( .A(net_12348), .Z(net_12349) );
XNOR2_X2 inst_326 ( .A(net_1026), .ZN(net_929), .B(net_192) );
SDFF_X2 inst_817 ( .SI(net_8508), .Q(net_8508), .D(net_3975), .SE(net_3884), .CK(net_12510) );
CLKBUF_X2 inst_10589 ( .A(net_10436), .Z(net_10437) );
CLKBUF_X2 inst_12550 ( .A(net_12397), .Z(net_12398) );
SDFFR_X2 inst_2194 ( .SI(net_6754), .Q(net_6754), .SE(net_2933), .D(net_2932), .CK(net_9111), .RN(x6501) );
CLKBUF_X2 inst_10789 ( .A(net_10636), .Z(net_10637) );
CLKBUF_X2 inst_16365 ( .A(net_16034), .Z(net_16213) );
CLKBUF_X2 inst_18419 ( .A(net_18266), .Z(net_18267) );
CLKBUF_X2 inst_18698 ( .A(net_18545), .Z(net_18546) );
CLKBUF_X2 inst_18691 ( .A(net_10508), .Z(net_18539) );
NOR3_X2 inst_3293 ( .A3(net_6157), .ZN(net_2167), .A2(net_2019), .A1(net_1350) );
CLKBUF_X2 inst_15825 ( .A(net_15672), .Z(net_15673) );
CLKBUF_X2 inst_18809 ( .A(net_18656), .Z(net_18657) );
CLKBUF_X2 inst_16808 ( .A(net_13377), .Z(net_16656) );
NAND4_X2 inst_3793 ( .ZN(net_3633), .A1(net_3516), .A2(net_3515), .A3(net_3514), .A4(net_3513) );
CLKBUF_X2 inst_18333 ( .A(net_14291), .Z(net_18181) );
XNOR2_X2 inst_108 ( .ZN(net_5467), .B(net_5019), .A(net_2117) );
CLKBUF_X2 inst_11143 ( .A(net_10990), .Z(net_10991) );
NAND2_X2 inst_4799 ( .ZN(net_1636), .A2(net_1376), .A1(net_726) );
NAND4_X2 inst_3778 ( .ZN(net_4243), .A1(net_3717), .A2(net_3716), .A3(net_3715), .A4(net_3714) );
CLKBUF_X2 inst_16475 ( .A(net_13103), .Z(net_16323) );
NAND3_X2 inst_3940 ( .ZN(net_4919), .A3(net_4678), .A1(net_4663), .A2(net_4643) );
INV_X2 inst_6503 ( .A(net_7584), .ZN(net_3107) );
SDFF_X2 inst_638 ( .SI(net_8553), .Q(net_8553), .SE(net_3979), .D(net_3939), .CK(net_12538) );
CLKBUF_X2 inst_11937 ( .A(net_11784), .Z(net_11785) );
AOI22_X2 inst_7786 ( .A1(net_5268), .B2(net_5267), .ZN(net_4864), .A2(net_4629), .B1(net_164) );
CLKBUF_X2 inst_10311 ( .A(net_10158), .Z(net_10159) );
CLKBUF_X2 inst_18139 ( .A(net_17817), .Z(net_17987) );
INV_X8 inst_5008 ( .ZN(net_4901), .A(net_4816) );
NOR3_X2 inst_3275 ( .A1(net_2415), .ZN(net_2411), .A3(net_2397), .A2(net_1776) );
CLKBUF_X2 inst_9237 ( .A(net_9084), .Z(net_9085) );
SDFF_X2 inst_1466 ( .SI(net_7291), .Q(net_7148), .D(net_7148), .SE(net_6279), .CK(net_17705) );
SDFF_X2 inst_1726 ( .Q(net_7993), .D(net_7993), .SI(net_2719), .SE(net_2542), .CK(net_15575) );
OR2_X4 inst_2841 ( .A2(net_2333), .ZN(net_2013), .A1(net_2012) );
DFFR_X2 inst_7157 ( .QN(net_7364), .D(net_2869), .CK(net_11836), .RN(x6501) );
CLKBUF_X2 inst_15591 ( .A(net_15438), .Z(net_15439) );
CLKBUF_X2 inst_14251 ( .A(net_10605), .Z(net_14099) );
DFFR_X2 inst_7118 ( .QN(net_7612), .D(net_3045), .CK(net_11926), .RN(x6501) );
CLKBUF_X2 inst_16170 ( .A(net_16017), .Z(net_16018) );
CLKBUF_X2 inst_10892 ( .A(net_10739), .Z(net_10740) );
CLKBUF_X2 inst_14576 ( .A(net_10812), .Z(net_14424) );
SDFF_X2 inst_905 ( .SI(net_8723), .Q(net_8723), .SE(net_6195), .D(net_3974), .CK(net_10814) );
CLKBUF_X2 inst_14677 ( .A(net_12343), .Z(net_14525) );
CLKBUF_X2 inst_16426 ( .A(net_13554), .Z(net_16274) );
CLKBUF_X2 inst_15991 ( .A(net_15838), .Z(net_15839) );
CLKBUF_X2 inst_11571 ( .A(net_9390), .Z(net_11419) );
CLKBUF_X2 inst_14860 ( .A(net_14707), .Z(net_14708) );
NAND2_X2 inst_4214 ( .A1(net_7011), .A2(net_5249), .ZN(net_5246) );
CLKBUF_X2 inst_12753 ( .A(net_12600), .Z(net_12601) );
CLKBUF_X2 inst_18242 ( .A(net_16403), .Z(net_18090) );
NAND4_X2 inst_3834 ( .ZN(net_2500), .A1(net_2344), .A4(net_2315), .A2(net_2163), .A3(net_2047) );
CLKBUF_X2 inst_16687 ( .A(net_16534), .Z(net_16535) );
NAND4_X2 inst_3651 ( .A4(net_6002), .A1(net_6001), .ZN(net_4614), .A2(net_4186), .A3(net_4185) );
SDFF_X2 inst_1759 ( .SI(net_7765), .Q(net_7765), .D(net_2639), .SE(net_2560), .CK(net_14388) );
SDFFR_X2 inst_2615 ( .Q(net_7366), .D(net_7366), .SE(net_1136), .CK(net_18640), .RN(x6501), .SI(x4861) );
CLKBUF_X2 inst_11792 ( .A(net_9752), .Z(net_11640) );
INV_X4 inst_5485 ( .A(net_1262), .ZN(net_861) );
CLKBUF_X2 inst_13859 ( .A(net_12680), .Z(net_13707) );
DFFR_X2 inst_7017 ( .QN(net_6290), .D(net_5729), .CK(net_13874), .RN(x6501) );
NOR2_X2 inst_3463 ( .ZN(net_2773), .A1(net_2438), .A2(net_2437) );
CLKBUF_X2 inst_16055 ( .A(net_15902), .Z(net_15903) );
CLKBUF_X2 inst_17867 ( .A(net_15288), .Z(net_17715) );
INV_X2 inst_6375 ( .A(net_3308), .ZN(net_1375) );
CLKBUF_X2 inst_11115 ( .A(net_10446), .Z(net_10963) );
CLKBUF_X2 inst_12492 ( .A(net_12339), .Z(net_12340) );
NAND2_X2 inst_4055 ( .ZN(net_5930), .A2(net_5927), .A1(net_2515) );
SDFF_X2 inst_1247 ( .SI(net_7691), .Q(net_7691), .SE(net_2714), .D(net_2713), .CK(net_14447) );
CLKBUF_X2 inst_16463 ( .A(net_15278), .Z(net_16311) );
INV_X4 inst_5284 ( .ZN(net_1769), .A(net_1621) );
CLKBUF_X2 inst_18942 ( .A(net_10168), .Z(net_18790) );
CLKBUF_X2 inst_13275 ( .A(net_13122), .Z(net_13123) );
CLKBUF_X2 inst_14541 ( .A(net_9446), .Z(net_14389) );
CLKBUF_X2 inst_17140 ( .A(net_16987), .Z(net_16988) );
SDFF_X2 inst_1493 ( .SI(net_7840), .Q(net_7840), .D(net_2721), .SE(net_2558), .CK(net_15773) );
OAI21_X2 inst_2998 ( .B2(net_5902), .ZN(net_5895), .A(net_5818), .B1(net_779) );
CLKBUF_X2 inst_11734 ( .A(net_11581), .Z(net_11582) );
SDFFR_X2 inst_2612 ( .Q(net_7386), .D(net_2803), .SE(net_1136), .CK(net_14954), .RN(x6501), .SI(x4607) );
CLKBUF_X2 inst_13348 ( .A(net_13195), .Z(net_13196) );
CLKBUF_X2 inst_14116 ( .A(net_13963), .Z(net_13964) );
CLKBUF_X2 inst_15623 ( .A(net_14350), .Z(net_15471) );
SDFF_X2 inst_1362 ( .Q(net_8200), .D(net_8200), .SI(net_2718), .SE(net_2561), .CK(net_14933) );
AOI21_X2 inst_8881 ( .ZN(net_5862), .A(net_5861), .B2(net_5784), .B1(x508) );
CLKBUF_X2 inst_12888 ( .A(net_12224), .Z(net_12736) );
CLKBUF_X2 inst_13798 ( .A(net_11482), .Z(net_13646) );
CLKBUF_X2 inst_19110 ( .A(net_17943), .Z(net_18958) );
XNOR2_X2 inst_272 ( .A(net_7582), .B(net_3990), .ZN(net_1041) );
CLKBUF_X2 inst_14311 ( .A(net_14158), .Z(net_14159) );
NAND2_X2 inst_4718 ( .A1(net_7371), .ZN(net_1972), .A2(net_1784) );
CLKBUF_X2 inst_9213 ( .A(net_9060), .Z(net_9061) );
NAND2_X2 inst_4133 ( .ZN(net_5389), .A1(net_5221), .A2(net_5003) );
SDFF_X2 inst_789 ( .SI(net_8360), .Q(net_8360), .D(net_3975), .SE(net_3880), .CK(net_12520) );
SDFF_X2 inst_1806 ( .D(net_7302), .SI(net_6959), .Q(net_6959), .SE(net_6281), .CK(net_18595) );
SDFF_X2 inst_1810 ( .SI(net_8059), .Q(net_8059), .D(net_2576), .SE(net_2508), .CK(net_15961) );
SDFF_X2 inst_1860 ( .D(net_7290), .SI(net_6947), .Q(net_6947), .SE(net_6281), .CK(net_15328) );
CLKBUF_X2 inst_15177 ( .A(net_15024), .Z(net_15025) );
CLKBUF_X2 inst_16636 ( .A(net_16483), .Z(net_16484) );
CLKBUF_X2 inst_15561 ( .A(net_15408), .Z(net_15409) );
SDFF_X2 inst_1885 ( .D(net_7296), .SI(net_6993), .Q(net_6993), .SE(net_6283), .CK(net_15811) );
CLKBUF_X2 inst_13232 ( .A(net_13079), .Z(net_13080) );
AOI22_X2 inst_7926 ( .A1(net_7942), .B1(net_7772), .A2(net_6092), .B2(net_6091), .ZN(net_4198) );
CLKBUF_X2 inst_11184 ( .A(net_11031), .Z(net_11032) );
CLKBUF_X2 inst_18505 ( .A(net_12424), .Z(net_18353) );
CLKBUF_X2 inst_14136 ( .A(net_13983), .Z(net_13984) );
CLKBUF_X2 inst_13189 ( .A(net_13036), .Z(net_13037) );
CLKBUF_X2 inst_18981 ( .A(net_18828), .Z(net_18829) );
NAND2_X2 inst_4885 ( .A2(net_7388), .ZN(net_712), .A1(net_177) );
CLKBUF_X2 inst_17149 ( .A(net_12605), .Z(net_16997) );
CLKBUF_X2 inst_18255 ( .A(net_18102), .Z(net_18103) );
SDFFR_X2 inst_2496 ( .Q(net_8980), .D(net_8980), .SI(net_4736), .SE(net_2562), .CK(net_16637), .RN(x6501) );
AOI22_X2 inst_8393 ( .B1(net_8747), .A1(net_8377), .A2(net_3867), .B2(net_3866), .ZN(net_3657) );
CLKBUF_X2 inst_13466 ( .A(net_13313), .Z(net_13314) );
CLKBUF_X2 inst_15158 ( .A(net_15005), .Z(net_15006) );
NAND2_X2 inst_4381 ( .A1(net_7117), .A2(net_5164), .ZN(net_5076) );
CLKBUF_X2 inst_17940 ( .A(net_17787), .Z(net_17788) );
CLKBUF_X2 inst_11406 ( .A(net_11253), .Z(net_11254) );
CLKBUF_X2 inst_11280 ( .A(net_9081), .Z(net_11128) );
AOI22_X2 inst_8229 ( .A1(net_8611), .B1(net_8426), .A2(net_3864), .B2(net_3863), .ZN(net_3808) );
SDFFR_X1 inst_2671 ( .D(net_6760), .SE(net_4506), .CK(net_11526), .RN(x6501), .SI(x2068), .Q(x2068) );
CLKBUF_X2 inst_17689 ( .A(net_17536), .Z(net_17537) );
CLKBUF_X2 inst_16675 ( .A(net_15076), .Z(net_16523) );
CLKBUF_X2 inst_9638 ( .A(net_9485), .Z(net_9486) );
CLKBUF_X2 inst_18118 ( .A(net_12009), .Z(net_17966) );
CLKBUF_X2 inst_14713 ( .A(net_13069), .Z(net_14561) );
CLKBUF_X2 inst_13068 ( .A(net_10416), .Z(net_12916) );
SDFF_X2 inst_1355 ( .Q(net_8199), .D(net_8199), .SI(net_2722), .SE(net_2561), .CK(net_14936) );
INV_X2 inst_6612 ( .A(net_7415), .ZN(net_6203) );
SDFF_X2 inst_877 ( .Q(net_8588), .D(net_8588), .SI(net_3950), .SE(net_3878), .CK(net_10962) );
CLKBUF_X2 inst_10267 ( .A(net_9807), .Z(net_10115) );
CLKBUF_X2 inst_18717 ( .A(net_18564), .Z(net_18565) );
INV_X2 inst_6563 ( .A(net_6807), .ZN(net_4622) );
CLKBUF_X2 inst_10704 ( .A(net_9847), .Z(net_10552) );
CLKBUF_X2 inst_12698 ( .A(net_12545), .Z(net_12546) );
DFFR_X1 inst_7372 ( .QN(net_5946), .D(net_5889), .CK(net_9410), .RN(x6501) );
INV_X2 inst_6384 ( .ZN(net_1329), .A(net_1328) );
CLKBUF_X2 inst_17430 ( .A(net_17277), .Z(net_17278) );
INV_X4 inst_5829 ( .A(net_7355), .ZN(net_1446) );
CLKBUF_X2 inst_14523 ( .A(net_14370), .Z(net_14371) );
INV_X4 inst_5904 ( .A(net_7484), .ZN(net_676) );
CLKBUF_X2 inst_10274 ( .A(net_9904), .Z(net_10122) );
CLKBUF_X2 inst_10734 ( .A(net_10581), .Z(net_10582) );
CLKBUF_X2 inst_11013 ( .A(net_10860), .Z(net_10861) );
AND2_X2 inst_9206 ( .ZN(net_1307), .A1(net_1188), .A2(net_883) );
SDFF_X2 inst_1894 ( .D(net_7277), .SI(net_6854), .Q(net_6854), .SE(net_6282), .CK(net_17347) );
CLKBUF_X2 inst_13960 ( .A(net_11967), .Z(net_13808) );
HA_X1 inst_6707 ( .S(net_2175), .CO(net_2088), .B(net_1604), .A(net_813) );
CLKBUF_X2 inst_15401 ( .A(net_15248), .Z(net_15249) );
NAND2_X2 inst_4643 ( .ZN(net_2445), .A2(net_2208), .A1(net_2008) );
CLKBUF_X2 inst_14379 ( .A(net_13547), .Z(net_14227) );
INV_X16 inst_6636 ( .ZN(net_3964), .A(net_3357) );
CLKBUF_X2 inst_13677 ( .A(net_13524), .Z(net_13525) );
SDFFR_X1 inst_2701 ( .SI(net_7533), .SE(net_5043), .CK(net_11934), .RN(x6501), .Q(x4143), .D(x4143) );
AOI22_X2 inst_8321 ( .B1(net_8808), .A1(net_8549), .A2(net_3861), .B2(net_3860), .ZN(net_3725) );
AND2_X2 inst_9171 ( .ZN(net_2753), .A1(net_2494), .A2(net_2383) );
CLKBUF_X2 inst_18078 ( .A(net_17925), .Z(net_17926) );
CLKBUF_X2 inst_10385 ( .A(net_10232), .Z(net_10233) );
OAI21_X2 inst_3165 ( .ZN(net_1651), .B1(net_1650), .A(net_1433), .B2(net_201) );
CLKBUF_X2 inst_11222 ( .A(net_11069), .Z(net_11070) );
SDFF_X2 inst_575 ( .Q(net_8840), .D(net_8840), .SE(net_3964), .SI(net_3954), .CK(net_12623) );
CLKBUF_X2 inst_11738 ( .A(net_11585), .Z(net_11586) );
CLKBUF_X2 inst_10151 ( .A(net_9998), .Z(net_9999) );
CLKBUF_X2 inst_16335 ( .A(net_14228), .Z(net_16183) );
CLKBUF_X2 inst_18130 ( .A(net_12998), .Z(net_17978) );
SDFF_X2 inst_627 ( .SI(net_8539), .Q(net_8539), .SE(net_3979), .D(net_3957), .CK(net_11009) );
CLKBUF_X2 inst_14606 ( .A(net_14453), .Z(net_14454) );
DFF_X1 inst_6831 ( .Q(net_6451), .D(net_3617), .CK(net_15169) );
NAND2_X2 inst_4725 ( .A1(net_7368), .ZN(net_1968), .A2(net_1783) );
NOR2_X2 inst_3352 ( .ZN(net_5573), .A1(net_5420), .A2(net_5419) );
SDFF_X2 inst_344 ( .SI(net_8481), .Q(net_8481), .SE(net_3983), .D(net_3948), .CK(net_13491) );
DFFS_X1 inst_6928 ( .D(net_6145), .CK(net_16362), .SN(x6501), .Q(x827) );
CLKBUF_X2 inst_17285 ( .A(net_17132), .Z(net_17133) );
NAND4_X2 inst_3818 ( .ZN(net_3608), .A1(net_3415), .A2(net_3414), .A3(net_3413), .A4(net_3412) );
INV_X4 inst_5975 ( .A(net_7498), .ZN(net_3544) );
CLKBUF_X2 inst_15209 ( .A(net_15056), .Z(net_15057) );
SDFF_X2 inst_1338 ( .Q(net_7949), .D(net_7949), .SE(net_2755), .SI(net_2658), .CK(net_18877) );
CLKBUF_X2 inst_17698 ( .A(net_17545), .Z(net_17546) );
SDFFR_X2 inst_2430 ( .SE(net_2678), .D(net_2512), .SI(net_444), .Q(net_444), .CK(net_13838), .RN(x6501) );
CLKBUF_X2 inst_13093 ( .A(net_9352), .Z(net_12941) );
MUX2_X2 inst_4952 ( .A(net_7382), .Z(net_2372), .S(net_2370), .B(net_815) );
NAND4_X2 inst_3731 ( .ZN(net_4299), .A1(net_4130), .A2(net_4129), .A3(net_4128), .A4(net_4127) );
CLKBUF_X2 inst_13932 ( .A(net_13779), .Z(net_13780) );
DFFS_X2 inst_6899 ( .Q(net_7481), .D(net_2524), .CK(net_16146), .SN(x6501) );
NAND2_X2 inst_4839 ( .A2(net_8890), .A1(net_3587), .ZN(net_1407) );
SDFF_X2 inst_2028 ( .SI(net_7917), .Q(net_7917), .D(net_2573), .SE(net_2461), .CK(net_15223) );
CLKBUF_X2 inst_15364 ( .A(net_12490), .Z(net_15212) );
AOI22_X2 inst_8381 ( .B1(net_8856), .A1(net_8301), .B2(net_6252), .A2(net_4345), .ZN(net_3667) );
CLKBUF_X2 inst_15038 ( .A(net_14885), .Z(net_14886) );
CLKBUF_X2 inst_16409 ( .A(net_16256), .Z(net_16257) );
CLKBUF_X2 inst_16994 ( .A(net_11080), .Z(net_16842) );
CLKBUF_X2 inst_14904 ( .A(net_14751), .Z(net_14752) );
SDFF_X2 inst_722 ( .SI(net_8490), .Q(net_8490), .D(net_3937), .SE(net_3884), .CK(net_10719) );
INV_X4 inst_6019 ( .ZN(net_2699), .A(net_162) );
AOI22_X2 inst_8093 ( .B1(net_8211), .A1(net_7701), .B2(net_6099), .A2(net_4399), .ZN(net_4054) );
CLKBUF_X2 inst_9502 ( .A(net_9323), .Z(net_9350) );
NAND2_X2 inst_4232 ( .A1(net_7001), .A2(net_5249), .ZN(net_5228) );
NAND2_X2 inst_4270 ( .A1(net_7037), .A2(net_5249), .ZN(net_5190) );
OAI21_X2 inst_3010 ( .B2(net_5755), .ZN(net_5720), .A(net_5719), .B1(net_720) );
CLKBUF_X2 inst_16726 ( .A(net_16573), .Z(net_16574) );
AOI22_X2 inst_8010 ( .B1(net_8132), .A1(net_7894), .A2(net_6098), .B2(net_4190), .ZN(net_4125) );
CLKBUF_X2 inst_17151 ( .A(net_16998), .Z(net_16999) );
CLKBUF_X2 inst_12282 ( .A(net_12129), .Z(net_12130) );
OAI21_X2 inst_3133 ( .B2(net_2204), .ZN(net_2103), .A(net_2102), .B1(net_2101) );
AOI22_X2 inst_8207 ( .B1(net_8682), .A1(net_8645), .B2(net_6109), .A2(net_3857), .ZN(net_3829) );
INV_X2 inst_6412 ( .A(net_6380), .ZN(net_871) );
SDFFR_X2 inst_2588 ( .Q(net_7297), .SI(net_7261), .D(net_1461), .SE(net_1327), .CK(net_15022), .RN(x6501) );
INV_X2 inst_6547 ( .A(net_7499), .ZN(net_510) );
CLKBUF_X2 inst_15844 ( .A(net_15691), .Z(net_15692) );
CLKBUF_X2 inst_15859 ( .A(net_10182), .Z(net_15707) );
CLKBUF_X2 inst_17671 ( .A(net_10617), .Z(net_17519) );
DFFR_X2 inst_6994 ( .QN(net_5977), .D(net_5870), .CK(net_10454), .RN(x6501) );
NAND2_X2 inst_4665 ( .ZN(net_2194), .A2(net_2005), .A1(net_1285) );
CLKBUF_X2 inst_15379 ( .A(net_15226), .Z(net_15227) );
CLKBUF_X2 inst_18142 ( .A(net_17989), .Z(net_17990) );
CLKBUF_X2 inst_18209 ( .A(net_12870), .Z(net_18057) );
CLKBUF_X2 inst_18837 ( .A(net_17272), .Z(net_18685) );
INV_X4 inst_5712 ( .A(net_7417), .ZN(net_609) );
INV_X4 inst_5562 ( .A(net_1854), .ZN(net_606) );
INV_X4 inst_5374 ( .A(net_1481), .ZN(net_1125) );
NAND2_X2 inst_4466 ( .A2(net_4783), .ZN(net_4781), .A1(x1152) );
CLKBUF_X2 inst_11058 ( .A(net_10534), .Z(net_10906) );
CLKBUF_X2 inst_15543 ( .A(net_9405), .Z(net_15391) );
CLKBUF_X2 inst_11035 ( .A(net_9582), .Z(net_10883) );
OR2_X2 inst_2875 ( .ZN(net_4395), .A1(net_4394), .A2(net_4393) );
AOI22_X2 inst_8447 ( .B1(net_6602), .A1(net_6569), .A2(net_6257), .B2(net_6110), .ZN(net_3493) );
AND2_X4 inst_9067 ( .ZN(net_3356), .A1(net_3245), .A2(net_3211) );
CLKBUF_X2 inst_11084 ( .A(net_10931), .Z(net_10932) );
CLKBUF_X2 inst_10341 ( .A(net_10188), .Z(net_10189) );
DFFR_X2 inst_7162 ( .QN(net_8902), .D(net_2780), .CK(net_16319), .RN(x6501) );
CLKBUF_X2 inst_9396 ( .A(net_9243), .Z(net_9244) );
INV_X2 inst_6248 ( .ZN(net_4858), .A(net_4752) );
NOR2_X2 inst_3389 ( .A2(net_4553), .ZN(net_4475), .A1(net_1605) );
SDFF_X2 inst_782 ( .SI(net_8351), .Q(net_8351), .D(net_3967), .SE(net_3880), .CK(net_10822) );
INV_X4 inst_5744 ( .A(net_7398), .ZN(net_726) );
OR2_X2 inst_2869 ( .ZN(net_5725), .A2(net_5712), .A1(net_5674) );
CLKBUF_X2 inst_10546 ( .A(net_10393), .Z(net_10394) );
XOR2_X2 inst_6 ( .Z(net_2885), .A(net_2565), .B(x3122) );
CLKBUF_X2 inst_10603 ( .A(net_10450), .Z(net_10451) );
CLKBUF_X2 inst_16181 ( .A(net_16028), .Z(net_16029) );
SDFFR_X2 inst_2486 ( .D(net_7368), .SE(net_2548), .SI(net_261), .Q(net_261), .CK(net_13546), .RN(x6501) );
INV_X4 inst_5461 ( .A(net_1856), .ZN(net_764) );
SDFFR_X2 inst_2410 ( .SE(net_2260), .Q(net_361), .D(net_361), .CK(net_9231), .RN(x6501), .SI(x1912) );
CLKBUF_X2 inst_11832 ( .A(net_11679), .Z(net_11680) );
AOI21_X2 inst_8927 ( .B2(net_5871), .ZN(net_5686), .A(net_5675), .B1(net_2684) );
AOI221_X4 inst_8728 ( .B1(net_8844), .C1(net_8363), .C2(net_6265), .B2(net_6253), .ZN(net_4337), .A(net_4246) );
CLKBUF_X2 inst_16670 ( .A(net_15634), .Z(net_16518) );
CLKBUF_X2 inst_12760 ( .A(net_11858), .Z(net_12608) );
CLKBUF_X2 inst_17674 ( .A(net_17521), .Z(net_17522) );
CLKBUF_X2 inst_14650 ( .A(net_14497), .Z(net_14498) );
CLKBUF_X2 inst_11726 ( .A(net_11573), .Z(net_11574) );
CLKBUF_X2 inst_17601 ( .A(net_17448), .Z(net_17449) );
CLKBUF_X2 inst_13030 ( .A(net_12877), .Z(net_12878) );
AOI22_X2 inst_8108 ( .B1(net_8145), .A1(net_7907), .A2(net_6098), .B2(net_4190), .ZN(net_4039) );
AOI22_X2 inst_8211 ( .A1(net_8609), .B1(net_8424), .A2(net_3864), .B2(net_3863), .ZN(net_3825) );
INV_X4 inst_6031 ( .A(net_8960), .ZN(net_1756) );
CLKBUF_X1 inst_7729 ( .A(x192486), .Z(x1016) );
SDFF_X2 inst_1026 ( .SI(net_7341), .Q(net_6748), .D(net_6748), .SE(net_3124), .CK(net_11901) );
SDFF_X2 inst_1320 ( .SI(net_7699), .Q(net_7699), .SE(net_2714), .D(net_2660), .CK(net_17021) );
CLKBUF_X2 inst_15638 ( .A(net_15485), .Z(net_15486) );
INV_X2 inst_6250 ( .ZN(net_4856), .A(net_4744) );
CLKBUF_X2 inst_11289 ( .A(net_10737), .Z(net_11137) );
INV_X4 inst_5576 ( .A(net_6393), .ZN(net_1949) );
CLKBUF_X2 inst_12826 ( .A(net_12673), .Z(net_12674) );
INV_X4 inst_5246 ( .A(net_2767), .ZN(net_2074) );
XOR2_X1 inst_95 ( .Z(net_1400), .B(net_1399), .A(net_775) );
NOR2_X2 inst_3376 ( .ZN(net_5549), .A2(net_5321), .A1(net_5320) );
OAI22_X2 inst_2921 ( .ZN(net_3209), .A2(net_3006), .B2(net_2537), .A1(net_1081), .B1(net_1080) );
CLKBUF_X2 inst_13058 ( .A(net_11448), .Z(net_12906) );
CLKBUF_X2 inst_10622 ( .A(net_10469), .Z(net_10470) );
CLKBUF_X2 inst_10499 ( .A(net_10346), .Z(net_10347) );
CLKBUF_X2 inst_14794 ( .A(net_11757), .Z(net_14642) );
CLKBUF_X2 inst_18358 ( .A(net_10605), .Z(net_18206) );
NAND3_X2 inst_4009 ( .ZN(net_1577), .A2(net_1083), .A3(net_827), .A1(net_502) );
CLKBUF_X2 inst_9766 ( .A(net_9613), .Z(net_9614) );
CLKBUF_X2 inst_10870 ( .A(net_10717), .Z(net_10718) );
AOI22_X2 inst_8071 ( .B1(net_8039), .A1(net_8005), .B2(net_6102), .A2(net_6097), .ZN(net_6046) );
AOI22_X2 inst_8297 ( .B1(net_8879), .A1(net_8324), .B2(net_6252), .A2(net_4345), .ZN(net_3745) );
NAND2_X2 inst_4900 ( .A2(net_7383), .ZN(net_620), .A1(net_172) );
CLKBUF_X2 inst_13325 ( .A(net_10042), .Z(net_13173) );
INV_X4 inst_5837 ( .A(net_7517), .ZN(net_538) );
INV_X4 inst_5394 ( .ZN(net_1054), .A(net_622) );
DFFR_X2 inst_7194 ( .QN(net_7161), .D(net_2434), .CK(net_18661), .RN(x6501) );
CLKBUF_X2 inst_13883 ( .A(net_13730), .Z(net_13731) );
DFFR_X1 inst_7537 ( .D(net_2696), .Q(net_293), .CK(net_11637), .RN(x6501) );
CLKBUF_X2 inst_17317 ( .A(net_17164), .Z(net_17165) );
CLKBUF_X2 inst_10407 ( .A(net_10254), .Z(net_10255) );
CLKBUF_X2 inst_19126 ( .A(net_16109), .Z(net_18974) );
CLKBUF_X2 inst_12369 ( .A(net_10765), .Z(net_12217) );
CLKBUF_X2 inst_19154 ( .A(net_19001), .Z(net_19002) );
AOI21_X2 inst_8955 ( .A(net_5746), .ZN(net_5602), .B1(net_5261), .B2(net_5255) );
NAND2_X2 inst_4901 ( .A2(net_7165), .A1(net_7164), .ZN(net_805) );
CLKBUF_X2 inst_14758 ( .A(net_12902), .Z(net_14606) );
NOR2_X2 inst_3590 ( .A1(net_2039), .ZN(net_910), .A2(net_909) );
CLKBUF_X2 inst_18783 ( .A(net_18630), .Z(net_18631) );
CLKBUF_X2 inst_18071 ( .A(net_13194), .Z(net_17919) );
CLKBUF_X2 inst_17594 ( .A(net_13420), .Z(net_17442) );
CLKBUF_X2 inst_18830 ( .A(net_10001), .Z(net_18678) );
AOI22_X2 inst_8145 ( .B1(net_8017), .A1(net_7983), .B2(net_6102), .A2(net_6097), .ZN(net_4006) );
CLKBUF_X2 inst_9252 ( .A(net_9099), .Z(net_9100) );
MUX2_X2 inst_4974 ( .A(net_9027), .Z(net_3945), .B(net_3194), .S(net_622) );
AOI22_X2 inst_8582 ( .B2(net_6319), .ZN(net_1790), .B1(net_1254), .A2(net_1253), .A1(x4367) );
CLKBUF_X2 inst_10836 ( .A(net_9607), .Z(net_10684) );
CLKBUF_X2 inst_18189 ( .A(net_18036), .Z(net_18037) );
SDFFR_X2 inst_2476 ( .Q(net_8992), .D(net_8992), .SI(net_4518), .SE(net_2562), .CK(net_16645), .RN(x6501) );
CLKBUF_X2 inst_16660 ( .A(net_10591), .Z(net_16508) );
CLKBUF_X2 inst_12078 ( .A(net_9777), .Z(net_11926) );
AOI22_X2 inst_8116 ( .B2(net_8081), .A1(net_7741), .B1(net_6108), .A2(net_6096), .ZN(net_4032) );
CLKBUF_X2 inst_18305 ( .A(net_18152), .Z(net_18153) );
NAND2_X2 inst_4502 ( .A2(net_4555), .ZN(net_4384), .A1(net_4383) );
CLKBUF_X2 inst_14258 ( .A(net_14105), .Z(net_14106) );
INV_X4 inst_5624 ( .A(net_8907), .ZN(net_5033) );
DFFR_X1 inst_7451 ( .QN(net_8934), .D(net_4748), .CK(net_14586), .RN(x6501) );
DFFR_X1 inst_7458 ( .QN(net_6422), .D(net_4726), .CK(net_9598), .RN(x6501) );
CLKBUF_X2 inst_14072 ( .A(net_13919), .Z(net_13920) );
SDFF_X2 inst_1036 ( .SI(net_7320), .Q(net_6694), .D(net_6694), .SE(net_3125), .CK(net_9864) );
CLKBUF_X2 inst_10094 ( .A(net_9941), .Z(net_9942) );
CLKBUF_X2 inst_10334 ( .A(net_10181), .Z(net_10182) );
AOI222_X1 inst_8653 ( .A2(net_6266), .C1(net_6204), .B2(net_4365), .C2(net_4364), .ZN(net_3913), .B1(net_1359), .A1(x13950) );
INV_X4 inst_5694 ( .A(net_6306), .ZN(net_2750) );
CLKBUF_X2 inst_14700 ( .A(net_13966), .Z(net_14548) );
CLKBUF_X2 inst_12141 ( .A(net_11988), .Z(net_11989) );
NAND2_X2 inst_4613 ( .A2(net_6144), .ZN(net_2615), .A1(net_2614) );
INV_X4 inst_5852 ( .A(net_7611), .ZN(net_1053) );
SDFFR_X2 inst_2376 ( .SE(net_2260), .Q(net_324), .D(net_324), .CK(net_11499), .RN(x6501), .SI(x2948) );
AOI22_X2 inst_7925 ( .B1(net_8078), .A1(net_7738), .B2(net_6108), .A2(net_6096), .ZN(net_4199) );
DFFR_X1 inst_7496 ( .QN(net_7615), .D(net_3061), .CK(net_9819), .RN(x6501) );
DFFR_X2 inst_7050 ( .QN(net_7504), .D(net_4841), .CK(net_17247), .RN(x6501) );
NAND2_X2 inst_4360 ( .A1(net_7110), .A2(net_5164), .ZN(net_5097) );
CLKBUF_X2 inst_19086 ( .A(net_18933), .Z(net_18934) );
SDFF_X2 inst_860 ( .Q(net_8568), .D(net_8568), .SI(net_3945), .SE(net_3878), .CK(net_13312) );
SDFF_X2 inst_563 ( .Q(net_8825), .D(net_8825), .SE(net_3964), .SI(net_3960), .CK(net_13136) );
CLKBUF_X2 inst_14074 ( .A(net_12244), .Z(net_13922) );
NAND3_X2 inst_3962 ( .ZN(net_6183), .A2(net_2946), .A1(net_2534), .A3(net_2486) );
SDFF_X2 inst_943 ( .SI(net_7325), .Q(net_6699), .D(net_6699), .SE(net_3125), .CK(net_9143) );
INV_X4 inst_5314 ( .ZN(net_1472), .A(net_1471) );
CLKBUF_X2 inst_15714 ( .A(net_13989), .Z(net_15562) );
CLKBUF_X2 inst_18979 ( .A(net_18826), .Z(net_18827) );
NAND2_X2 inst_4711 ( .ZN(net_2025), .A1(net_1836), .A2(net_1835) );
SDFF_X2 inst_1964 ( .D(net_7288), .SI(net_7025), .Q(net_7025), .SE(net_6277), .CK(net_17661) );
CLKBUF_X2 inst_12151 ( .A(net_10302), .Z(net_11999) );
DFFR_X1 inst_7464 ( .QN(net_7440), .D(net_4377), .CK(net_12937), .RN(x6501) );
SDFF_X2 inst_1765 ( .SI(net_8070), .Q(net_8070), .D(net_2710), .SE(net_2508), .CK(net_14387) );
CLKBUF_X2 inst_18908 ( .A(net_13660), .Z(net_18756) );
CLKBUF_X2 inst_18657 ( .A(net_18504), .Z(net_18505) );
CLKBUF_X2 inst_13525 ( .A(net_12160), .Z(net_13373) );
INV_X2 inst_6357 ( .ZN(net_2195), .A(net_2105) );
CLKBUF_X2 inst_11944 ( .A(net_11791), .Z(net_11792) );
CLKBUF_X2 inst_17279 ( .A(net_17126), .Z(net_17127) );
CLKBUF_X2 inst_16231 ( .A(net_16078), .Z(net_16079) );
XNOR2_X2 inst_178 ( .ZN(net_1717), .A(net_1360), .B(net_938) );
CLKBUF_X2 inst_18588 ( .A(net_14253), .Z(net_18436) );
AND2_X2 inst_9179 ( .ZN(net_2231), .A1(net_2141), .A2(net_2140) );
AOI22_X2 inst_8257 ( .A1(net_8615), .B1(net_8430), .A2(net_3864), .B2(net_3863), .ZN(net_3781) );
INV_X4 inst_5941 ( .A(net_7243), .ZN(net_1961) );
CLKBUF_X2 inst_13562 ( .A(net_13082), .Z(net_13410) );
SDFF_X2 inst_1148 ( .SI(net_7329), .Q(net_6604), .D(net_6604), .SE(net_3069), .CK(net_11646) );
NAND3_X2 inst_3919 ( .ZN(net_5619), .A1(net_5548), .A3(net_5482), .A2(net_5315) );
CLKBUF_X2 inst_17643 ( .A(net_17490), .Z(net_17491) );
CLKBUF_X2 inst_10292 ( .A(net_10139), .Z(net_10140) );
NAND2_X2 inst_4350 ( .A1(net_7148), .A2(net_5166), .ZN(net_5107) );
AOI22_X2 inst_8270 ( .B1(net_8802), .A1(net_8543), .ZN(net_6226), .A2(net_3861), .B2(net_3860) );
CLKBUF_X2 inst_18467 ( .A(net_12324), .Z(net_18315) );
CLKBUF_X2 inst_9659 ( .A(net_9333), .Z(net_9507) );
INV_X4 inst_6004 ( .A(net_6304), .ZN(net_719) );
SDFF_X2 inst_842 ( .SI(net_8653), .Q(net_8653), .D(net_3942), .SE(net_3885), .CK(net_10511) );
SDFFS_X2 inst_2068 ( .SI(net_7390), .SE(net_2417), .Q(net_179), .D(net_179), .CK(net_14733), .SN(x6501) );
CLKBUF_X2 inst_9897 ( .A(net_9744), .Z(net_9745) );
SDFF_X2 inst_551 ( .Q(net_8669), .D(net_8669), .SI(net_3980), .SE(net_3935), .CK(net_13346) );
CLKBUF_X2 inst_9697 ( .A(net_9544), .Z(net_9545) );
CLKBUF_X2 inst_17577 ( .A(net_17424), .Z(net_17425) );
SDFFS_X1 inst_2101 ( .Q(net_6800), .D(net_6800), .SE(net_6272), .SI(net_1666), .CK(net_9537), .SN(x6501) );
SDFF_X2 inst_353 ( .Q(net_8748), .D(net_8748), .SE(net_3982), .SI(net_3981), .CK(net_10749) );
CLKBUF_X2 inst_19132 ( .A(net_12677), .Z(net_18980) );
NAND4_X2 inst_3808 ( .ZN(net_3618), .A1(net_3455), .A2(net_3454), .A3(net_3453), .A4(net_3452) );
CLKBUF_X2 inst_15721 ( .A(net_11569), .Z(net_15569) );
CLKBUF_X2 inst_18819 ( .A(net_10783), .Z(net_18667) );
SDFF_X2 inst_1940 ( .SI(net_8046), .Q(net_8046), .D(net_2705), .SE(net_2508), .CK(net_18519) );
INV_X2 inst_6286 ( .ZN(net_4214), .A(net_3923) );
CLKBUF_X2 inst_16770 ( .A(net_16617), .Z(net_16618) );
NAND2_X2 inst_4632 ( .A2(net_5871), .ZN(net_2513), .A1(net_2512) );
AOI22_X2 inst_8492 ( .B1(net_6546), .A1(net_6513), .A2(net_6137), .B2(net_6104), .ZN(net_3448) );
CLKBUF_X2 inst_10400 ( .A(net_10198), .Z(net_10248) );
CLKBUF_X2 inst_13456 ( .A(net_12012), .Z(net_13304) );
CLKBUF_X2 inst_15025 ( .A(net_14872), .Z(net_14873) );
INV_X2 inst_6212 ( .ZN(net_5498), .A(net_5381) );
CLKBUF_X2 inst_13917 ( .A(net_13764), .Z(net_13765) );
NAND2_X4 inst_4041 ( .A2(net_6276), .ZN(net_2474), .A1(net_2239) );
CLKBUF_X2 inst_13761 ( .A(net_13608), .Z(net_13609) );
CLKBUF_X2 inst_9559 ( .A(net_9406), .Z(net_9407) );
CLKBUF_X2 inst_14184 ( .A(net_14031), .Z(net_14032) );
CLKBUF_X2 inst_13869 ( .A(net_13716), .Z(net_13717) );
CLKBUF_X2 inst_14588 ( .A(net_14435), .Z(net_14436) );
DFF_X1 inst_6745 ( .QN(net_6789), .D(net_5624), .CK(net_9397) );
CLKBUF_X2 inst_11321 ( .A(net_11168), .Z(net_11169) );
CLKBUF_X2 inst_14064 ( .A(net_13911), .Z(net_13912) );
CLKBUF_X2 inst_18824 ( .A(net_18671), .Z(net_18672) );
CLKBUF_X2 inst_17626 ( .A(net_17473), .Z(net_17474) );
CLKBUF_X2 inst_13980 ( .A(net_11436), .Z(net_13828) );
CLKBUF_X2 inst_12624 ( .A(net_11395), .Z(net_12472) );
DFFR_X2 inst_7134 ( .QN(net_8949), .D(net_3025), .CK(net_17241), .RN(x6501) );
NOR2_X2 inst_3370 ( .ZN(net_5555), .A1(net_5348), .A2(net_5347) );
CLKBUF_X2 inst_10168 ( .A(net_9408), .Z(net_10016) );
CLKBUF_X2 inst_15301 ( .A(net_15148), .Z(net_15149) );
AOI21_X2 inst_8993 ( .B2(net_1779), .ZN(net_1438), .A(net_1034), .B1(net_205) );
INV_X2 inst_6579 ( .A(net_8902), .ZN(net_484) );
DFFR_X2 inst_7210 ( .D(net_2358), .QN(net_222), .CK(net_17565), .RN(x6501) );
SDFF_X2 inst_901 ( .SI(net_8718), .Q(net_8718), .SE(net_6195), .D(net_3959), .CK(net_9978) );
CLKBUF_X2 inst_10992 ( .A(net_10839), .Z(net_10840) );
DFFR_X2 inst_7261 ( .QN(net_7401), .D(net_1973), .CK(net_17860), .RN(x6501) );
INV_X4 inst_6094 ( .A(net_8913), .ZN(net_2622) );
CLKBUF_X2 inst_13821 ( .A(net_9998), .Z(net_13669) );
CLKBUF_X2 inst_9957 ( .A(net_9804), .Z(net_9805) );
CLKBUF_X2 inst_10863 ( .A(net_10710), .Z(net_10711) );
CLKBUF_X2 inst_14843 ( .A(net_13550), .Z(net_14691) );
SDFFR_X2 inst_2403 ( .SI(net_7379), .SE(net_2723), .D(net_2694), .QN(net_160), .CK(net_15036), .RN(x6501) );
MUX2_X2 inst_4948 ( .A(net_7375), .Z(net_2377), .S(net_2376), .B(net_889) );
AND2_X4 inst_9104 ( .A2(net_2299), .ZN(net_2268), .A1(net_1456) );
CLKBUF_X2 inst_14545 ( .A(net_14392), .Z(net_14393) );
OAI21_X2 inst_3098 ( .A(net_2892), .ZN(net_2769), .B1(net_2768), .B2(net_2767) );
CLKBUF_X2 inst_13834 ( .A(net_13681), .Z(net_13682) );
CLKBUF_X2 inst_10679 ( .A(net_10149), .Z(net_10527) );
INV_X4 inst_6144 ( .A(net_6134), .ZN(net_6133) );
INV_X8 inst_5013 ( .ZN(net_4898), .A(net_4396) );
CLKBUF_X2 inst_12034 ( .A(net_11881), .Z(net_11882) );
INV_X4 inst_5910 ( .A(net_7232), .ZN(net_1809) );
SDFF_X2 inst_928 ( .SI(net_8721), .Q(net_8721), .SE(net_6195), .D(net_3967), .CK(net_13078) );
CLKBUF_X2 inst_15782 ( .A(net_10508), .Z(net_15630) );
CLKBUF_X2 inst_10695 ( .A(net_10542), .Z(net_10543) );
CLKBUF_X2 inst_17828 ( .A(net_17675), .Z(net_17676) );
SDFF_X2 inst_1539 ( .Q(net_7992), .D(net_7992), .SI(net_2575), .SE(net_2542), .CK(net_15996) );
SDFFR_X1 inst_2662 ( .D(net_6784), .SE(net_4506), .CK(net_9181), .RN(x6501), .SI(x1305), .Q(x1305) );
CLKBUF_X2 inst_16309 ( .A(net_16156), .Z(net_16157) );
CLKBUF_X2 inst_18035 ( .A(net_17882), .Z(net_17883) );
SDFF_X2 inst_1718 ( .Q(net_8141), .D(net_8141), .SI(net_2660), .SE(net_2541), .CK(net_14252) );
CLKBUF_X2 inst_18912 ( .A(net_18759), .Z(net_18760) );
CLKBUF_X2 inst_9424 ( .A(net_9271), .Z(net_9272) );
AOI22_X2 inst_8549 ( .B2(net_4889), .A1(net_4803), .ZN(net_3389), .B1(net_3388), .A2(net_3238) );
CLKBUF_X2 inst_18385 ( .A(net_18232), .Z(net_18233) );
CLKBUF_X2 inst_11126 ( .A(net_10973), .Z(net_10974) );
CLKBUF_X2 inst_16779 ( .A(net_16626), .Z(net_16627) );
SDFF_X2 inst_1296 ( .Q(net_8098), .D(net_8098), .SI(net_2718), .SE(net_2707), .CK(net_18812) );
CLKBUF_X2 inst_14443 ( .A(net_9102), .Z(net_14291) );
NAND4_X2 inst_3671 ( .A4(net_6048), .A1(net_6047), .ZN(net_4594), .A2(net_4066), .A3(net_4065) );
CLKBUF_X2 inst_17781 ( .A(net_17628), .Z(net_17629) );
AOI22_X2 inst_7978 ( .B1(net_8026), .A1(net_7992), .B2(net_6102), .A2(net_6097), .ZN(net_4152) );
CLKBUF_X2 inst_13121 ( .A(net_12968), .Z(net_12969) );
NAND2_X2 inst_4513 ( .A2(net_6207), .A1(net_4320), .ZN(net_4318) );
CLKBUF_X2 inst_15078 ( .A(net_10762), .Z(net_14926) );
INV_X2 inst_6290 ( .ZN(net_4209), .A(net_3917) );
CLKBUF_X2 inst_10855 ( .A(net_10702), .Z(net_10703) );
CLKBUF_X2 inst_17339 ( .A(net_12664), .Z(net_17187) );
NAND2_X2 inst_4452 ( .ZN(net_4964), .A2(net_4962), .A1(net_3255) );
CLKBUF_X2 inst_10633 ( .A(net_10480), .Z(net_10481) );
CLKBUF_X2 inst_9954 ( .A(net_9801), .Z(net_9802) );
NAND2_X2 inst_4151 ( .ZN(net_5365), .A1(net_5209), .A2(net_4997) );
SDFF_X2 inst_1825 ( .D(net_7274), .SI(net_6851), .Q(net_6851), .SE(net_6282), .CK(net_14120) );
SDFF_X2 inst_1606 ( .Q(net_8142), .D(net_8142), .SI(net_2704), .SE(net_2541), .CK(net_14270) );
OR2_X4 inst_2851 ( .A1(net_7206), .ZN(net_1722), .A2(net_1374) );
INV_X4 inst_5619 ( .A(net_8955), .ZN(net_909) );
INV_X4 inst_5126 ( .ZN(net_4809), .A(net_4381) );
SDFF_X2 inst_410 ( .SI(net_8324), .Q(net_8324), .SE(net_3978), .D(net_3941), .CK(net_12909) );
XNOR2_X2 inst_316 ( .B(net_7396), .ZN(net_949), .A(net_948) );
SDFF_X2 inst_1174 ( .D(net_7326), .SI(net_6502), .Q(net_6502), .SE(net_3071), .CK(net_11275) );
CLKBUF_X2 inst_12860 ( .A(net_12707), .Z(net_12708) );
SDFF_X2 inst_1023 ( .SI(net_7319), .Q(net_6726), .D(net_6726), .SE(net_3124), .CK(net_12019) );
CLKBUF_X2 inst_16665 ( .A(net_10939), .Z(net_16513) );
CLKBUF_X2 inst_17509 ( .A(net_17356), .Z(net_17357) );
SDFF_X2 inst_678 ( .SI(net_8613), .Q(net_8613), .SE(net_3984), .D(net_3957), .CK(net_13251) );
AOI22_X2 inst_8515 ( .B1(net_6617), .A1(net_6584), .A2(net_6257), .B2(net_6110), .ZN(net_3425) );
CLKBUF_X2 inst_17429 ( .A(net_11284), .Z(net_17277) );
NAND2_X2 inst_4359 ( .A1(net_7150), .A2(net_5166), .ZN(net_5098) );
CLKBUF_X2 inst_16936 ( .A(net_16783), .Z(net_16784) );
DFFR_X2 inst_7310 ( .D(net_291), .QN(net_150), .CK(net_11141), .RN(x6501) );
CLKBUF_X2 inst_13177 ( .A(net_13024), .Z(net_13025) );
CLKBUF_X2 inst_15765 ( .A(net_15612), .Z(net_15613) );
AOI22_X2 inst_8033 ( .B1(net_7931), .A1(net_7829), .B2(net_6103), .A2(net_4398), .ZN(net_4105) );
CLKBUF_X2 inst_12191 ( .A(net_9313), .Z(net_12039) );
SDFF_X2 inst_1946 ( .SI(net_8050), .Q(net_8050), .D(net_2708), .SE(net_2508), .CK(net_18263) );
CLKBUF_X2 inst_10472 ( .A(net_10319), .Z(net_10320) );
AOI222_X1 inst_8686 ( .B1(net_6485), .A2(net_3296), .B2(net_3295), .C2(net_3294), .ZN(net_3285), .C1(net_3284), .A1(net_1214) );
INV_X4 inst_5322 ( .A(net_2424), .ZN(net_2244) );
CLKBUF_X2 inst_9226 ( .A(net_9064), .Z(net_9074) );
CLKBUF_X2 inst_9786 ( .A(net_9633), .Z(net_9634) );
AND2_X4 inst_9073 ( .ZN(net_6255), .A2(net_6082), .A1(net_6081) );
NOR2_X2 inst_3457 ( .ZN(net_2899), .A2(net_2850), .A1(net_2527) );
CLKBUF_X2 inst_12996 ( .A(net_12843), .Z(net_12844) );
SDFF_X2 inst_688 ( .Q(net_8861), .D(net_8861), .SI(net_3946), .SE(net_3936), .CK(net_11068) );
SDFFR_X2 inst_2549 ( .QN(net_6372), .SE(net_2147), .D(net_2135), .SI(net_1944), .CK(net_18138), .RN(x6501) );
NAND4_X2 inst_3641 ( .ZN(net_4943), .A1(net_4721), .A4(net_4579), .A3(net_4545), .A2(net_4482) );
NAND2_X2 inst_4894 ( .A2(net_7380), .ZN(net_651), .A1(net_169) );
SDFFR_X2 inst_2387 ( .SE(net_2260), .Q(net_375), .D(net_375), .CK(net_11392), .RN(x6501), .SI(x1500) );
CLKBUF_X2 inst_15372 ( .A(net_14472), .Z(net_15220) );
CLKBUF_X2 inst_16099 ( .A(net_15946), .Z(net_15947) );
CLKBUF_X2 inst_12980 ( .A(net_12827), .Z(net_12828) );
CLKBUF_X2 inst_13351 ( .A(net_10388), .Z(net_13199) );
CLKBUF_X2 inst_14416 ( .A(net_14263), .Z(net_14264) );
NAND2_X2 inst_4391 ( .A1(net_7043), .A2(net_5162), .ZN(net_5066) );
CLKBUF_X2 inst_12474 ( .A(net_12150), .Z(net_12322) );
CLKBUF_X2 inst_10137 ( .A(net_9795), .Z(net_9985) );
CLKBUF_X2 inst_10017 ( .A(net_9736), .Z(net_9865) );
CLKBUF_X2 inst_10163 ( .A(net_10010), .Z(net_10011) );
INV_X2 inst_6423 ( .ZN(net_750), .A(net_749) );
OAI21_X2 inst_3156 ( .B2(net_1984), .ZN(net_1975), .A(net_1974), .B1(net_1521) );
SDFFR_X1 inst_2747 ( .SI(net_9016), .Q(net_9016), .D(net_7445), .SE(net_3208), .CK(net_12830), .RN(x6501) );
CLKBUF_X2 inst_13744 ( .A(net_12738), .Z(net_13592) );
SDFF_X2 inst_1220 ( .Q(net_7955), .D(net_7955), .SE(net_2755), .SI(net_2720), .CK(net_18424) );
SDFF_X2 inst_1456 ( .SI(net_7273), .Q(net_7130), .D(net_7130), .SE(net_6279), .CK(net_14136) );
SDFFR_X2 inst_2181 ( .QN(net_7575), .D(net_3959), .SE(net_3144), .SI(net_3052), .CK(net_10871), .RN(x6501) );
AOI22_X2 inst_8554 ( .A2(net_6182), .B1(net_3161), .ZN(net_3002), .A1(net_1637), .B2(net_1302) );
AOI21_X2 inst_8909 ( .ZN(net_5788), .A(net_5745), .B2(net_5653), .B1(net_4935) );
CLKBUF_X2 inst_16904 ( .A(net_12480), .Z(net_16752) );
AOI21_X2 inst_8965 ( .ZN(net_3152), .B2(net_3072), .B1(net_2948), .A(net_2310) );
INV_X4 inst_5154 ( .ZN(net_3246), .A(net_3217) );
NAND2_X2 inst_4195 ( .ZN(net_5304), .A2(net_5180), .A1(net_5060) );
CLKBUF_X2 inst_10593 ( .A(net_10303), .Z(net_10441) );
AOI22_X2 inst_8473 ( .B1(net_6740), .A1(net_6707), .B2(net_6202), .A2(net_3520), .ZN(net_3467) );
CLKBUF_X2 inst_9305 ( .A(net_9152), .Z(net_9153) );
CLKBUF_X2 inst_13605 ( .A(net_13452), .Z(net_13453) );
NAND2_X2 inst_4440 ( .A1(net_6877), .A2(net_5016), .ZN(net_4987) );
DFFR_X2 inst_7072 ( .QN(net_8897), .D(net_4226), .CK(net_13534), .RN(x6501) );
INV_X4 inst_5959 ( .A(net_7435), .ZN(net_3274) );
CLKBUF_X2 inst_11607 ( .A(net_11297), .Z(net_11455) );
CLKBUF_X2 inst_17292 ( .A(net_14043), .Z(net_17140) );
AND2_X4 inst_9149 ( .ZN(net_6278), .A2(net_2265), .A1(net_1176) );
NAND2_X2 inst_4199 ( .ZN(net_5298), .A1(net_5177), .A2(net_4981) );
CLKBUF_X2 inst_18174 ( .A(net_18021), .Z(net_18022) );
CLKBUF_X2 inst_13588 ( .A(net_11902), .Z(net_13436) );
CLKBUF_X2 inst_14370 ( .A(net_9251), .Z(net_14218) );
CLKBUF_X2 inst_12718 ( .A(net_12565), .Z(net_12566) );
AOI21_X2 inst_8902 ( .ZN(net_5844), .A(net_5783), .B2(net_5690), .B1(net_4909) );
INV_X4 inst_5749 ( .A(net_7221), .ZN(net_1499) );
INV_X2 inst_6225 ( .ZN(net_5485), .A(net_5326) );
CLKBUF_X2 inst_12754 ( .A(net_12601), .Z(net_12602) );
NAND2_X2 inst_4420 ( .A1(net_6859), .A2(net_5016), .ZN(net_5007) );
CLKBUF_X2 inst_14209 ( .A(net_10897), .Z(net_14057) );
CLKBUF_X2 inst_13795 ( .A(net_13642), .Z(net_13643) );
SDFF_X2 inst_1057 ( .D(net_7314), .SI(net_6622), .Q(net_6622), .SE(net_3123), .CK(net_9933) );
CLKBUF_X2 inst_14097 ( .A(net_13944), .Z(net_13945) );
CLKBUF_X2 inst_10359 ( .A(net_10206), .Z(net_10207) );
CLKBUF_X2 inst_15225 ( .A(net_11093), .Z(net_15073) );
AOI221_X2 inst_8843 ( .B1(net_8051), .C1(net_7847), .B2(net_6107), .ZN(net_6031), .C2(net_4400), .A(net_4279) );
CLKBUF_X2 inst_17118 ( .A(net_16965), .Z(net_16966) );
INV_X4 inst_5191 ( .ZN(net_2967), .A(net_2943) );
CLKBUF_X2 inst_14565 ( .A(net_14412), .Z(net_14413) );
INV_X4 inst_5602 ( .A(net_7567), .ZN(net_593) );
CLKBUF_X2 inst_16497 ( .A(net_16344), .Z(net_16345) );
CLKBUF_X2 inst_10743 ( .A(net_10590), .Z(net_10591) );
CLKBUF_X2 inst_17487 ( .A(net_17334), .Z(net_17335) );
SDFF_X2 inst_748 ( .Q(net_8778), .D(net_8778), .SI(net_3961), .SE(net_3879), .CK(net_13182) );
CLKBUF_X2 inst_10610 ( .A(net_9287), .Z(net_10458) );
OR2_X4 inst_2839 ( .ZN(net_2225), .A1(net_2224), .A2(net_2223) );
AOI222_X1 inst_8609 ( .B2(net_6765), .B1(net_5835), .A2(net_5830), .C2(net_5824), .ZN(net_5804), .A1(net_2920), .C1(net_2132) );
DFF_X1 inst_6730 ( .Q(net_6775), .D(net_5639), .CK(net_9211) );
CLKBUF_X2 inst_17097 ( .A(net_16944), .Z(net_16945) );
CLKBUF_X2 inst_11373 ( .A(net_11015), .Z(net_11221) );
NAND2_X2 inst_4582 ( .A1(net_6459), .A2(net_3033), .ZN(net_2951) );
CLKBUF_X2 inst_9266 ( .A(net_9113), .Z(net_9114) );
CLKBUF_X2 inst_16973 ( .A(net_9406), .Z(net_16821) );
CLKBUF_X2 inst_18152 ( .A(net_11452), .Z(net_18000) );
INV_X4 inst_5532 ( .ZN(net_820), .A(net_658) );
NAND2_X2 inst_4526 ( .A2(net_3574), .ZN(net_3560), .A1(net_3557) );
CLKBUF_X2 inst_15700 ( .A(net_15547), .Z(net_15548) );
CLKBUF_X2 inst_11070 ( .A(net_10917), .Z(net_10918) );
CLKBUF_X2 inst_17406 ( .A(net_17253), .Z(net_17254) );
NAND2_X2 inst_4587 ( .ZN(net_2886), .A2(net_2763), .A1(net_1281) );
SDFF_X2 inst_1986 ( .D(net_7281), .SI(net_6898), .Q(net_6898), .SE(net_6284), .CK(net_18973) );
SDFF_X2 inst_1949 ( .D(net_7281), .SI(net_6938), .Q(net_6938), .SE(net_6281), .CK(net_18985) );
INV_X32 inst_6170 ( .ZN(net_5249), .A(net_4814) );
INV_X4 inst_5726 ( .A(net_7256), .ZN(net_1939) );
CLKBUF_X2 inst_10644 ( .A(net_10491), .Z(net_10492) );
CLKBUF_X2 inst_12163 ( .A(net_10005), .Z(net_12011) );
CLKBUF_X2 inst_15899 ( .A(net_9757), .Z(net_15747) );
INV_X4 inst_5867 ( .A(net_8928), .ZN(net_2606) );
AOI22_X2 inst_8243 ( .B1(net_8853), .A1(net_8298), .B2(net_6252), .A2(net_4345), .ZN(net_3794) );
OAI22_X2 inst_2911 ( .A2(net_8233), .B2(net_6133), .A1(net_4954), .ZN(net_4873), .B1(net_1509) );
CLKBUF_X2 inst_13770 ( .A(net_13617), .Z(net_13618) );
SDFF_X2 inst_1859 ( .D(net_7289), .SI(net_6946), .Q(net_6946), .SE(net_6281), .CK(net_15333) );
AOI22_X4 inst_7734 ( .A1(net_7974), .B1(net_7804), .A2(net_6092), .B2(net_6091), .ZN(net_4043) );
AOI22_X2 inst_8238 ( .A1(net_8594), .B1(net_8409), .A2(net_3864), .B2(net_3863), .ZN(net_3799) );
OR2_X4 inst_2815 ( .A1(net_7645), .A2(net_7644), .ZN(net_5272) );
CLKBUF_X2 inst_15818 ( .A(net_15665), .Z(net_15666) );
AOI22_X2 inst_8267 ( .B1(net_8579), .A1(net_8468), .A2(net_6263), .B2(net_6262), .ZN(net_3771) );
INV_X4 inst_5754 ( .A(net_7393), .ZN(net_1780) );
NAND2_X2 inst_4208 ( .ZN(net_5286), .A1(net_5171), .A2(net_4978) );
AOI22_X2 inst_8426 ( .B1(net_6663), .A1(net_6630), .A2(net_6213), .B2(net_6138), .ZN(net_3515) );
NOR2_X2 inst_3605 ( .ZN(net_824), .A1(net_560), .A2(net_269) );
SDFF_X2 inst_651 ( .Q(net_8423), .D(net_8423), .SI(net_3973), .SE(net_3934), .CK(net_10920) );
CLKBUF_X2 inst_9617 ( .A(net_9301), .Z(net_9465) );
CLKBUF_X2 inst_15977 ( .A(net_15824), .Z(net_15825) );
CLKBUF_X2 inst_11392 ( .A(net_11239), .Z(net_11240) );
SDFF_X2 inst_1157 ( .SI(net_7340), .Q(net_6615), .D(net_6615), .SE(net_3069), .CK(net_9607) );
CLKBUF_X2 inst_11560 ( .A(net_10842), .Z(net_11408) );
AOI22_X2 inst_8065 ( .A1(net_7970), .B1(net_7800), .A2(net_6092), .B2(net_6091), .ZN(net_4078) );
CLKBUF_X2 inst_9993 ( .A(net_9633), .Z(net_9841) );
AOI22_X2 inst_8408 ( .B1(net_8675), .A1(net_8638), .B2(net_6109), .A2(net_3857), .ZN(net_3644) );
CLKBUF_X2 inst_13395 ( .A(net_12237), .Z(net_13243) );
CLKBUF_X2 inst_16414 ( .A(net_15638), .Z(net_16262) );
NOR2_X2 inst_3528 ( .A1(net_1700), .ZN(net_1692), .A2(net_1113) );
SDFFS_X2 inst_2061 ( .Q(net_8271), .D(net_8271), .SI(net_6148), .SE(net_2996), .CK(net_18427), .SN(x6501) );
NAND2_X2 inst_4255 ( .A1(net_6882), .A2(net_5247), .ZN(net_5205) );
CLKBUF_X2 inst_13486 ( .A(net_12906), .Z(net_13334) );
INV_X4 inst_6138 ( .A(net_6120), .ZN(net_6115) );
CLKBUF_X2 inst_14981 ( .A(net_14821), .Z(net_14829) );
INV_X4 inst_5272 ( .ZN(net_1690), .A(net_1689) );
CLKBUF_X2 inst_15242 ( .A(net_14261), .Z(net_15090) );
CLKBUF_X2 inst_17980 ( .A(net_17827), .Z(net_17828) );
SDFFR_X2 inst_2262 ( .D(net_7379), .SE(net_2802), .SI(net_188), .Q(net_188), .CK(net_14976), .RN(x6501) );
NOR3_X2 inst_3288 ( .ZN(net_2256), .A2(net_2255), .A1(net_2083), .A3(net_1327) );
CLKBUF_X2 inst_18898 ( .A(net_18745), .Z(net_18746) );
SDFF_X2 inst_1160 ( .SI(net_7310), .Q(net_6618), .D(net_6618), .SE(net_3069), .CK(net_9605) );
SDFF_X2 inst_1394 ( .SI(net_7729), .Q(net_7729), .D(net_2711), .SE(net_2559), .CK(net_14289) );
AND2_X4 inst_9131 ( .ZN(net_1399), .A2(net_849), .A1(net_182) );
CLKBUF_X2 inst_13724 ( .A(net_13571), .Z(net_13572) );
CLKBUF_X2 inst_17951 ( .A(net_15966), .Z(net_17799) );
CLKBUF_X2 inst_10767 ( .A(net_10614), .Z(net_10615) );
SDFF_X2 inst_1876 ( .D(net_7264), .SI(net_6961), .Q(net_6961), .SE(net_6283), .CK(net_17415) );
CLKBUF_X2 inst_18517 ( .A(net_18364), .Z(net_18365) );
CLKBUF_X2 inst_12869 ( .A(net_12716), .Z(net_12717) );
SDFF_X2 inst_1315 ( .SI(net_7702), .Q(net_7702), .SE(net_2714), .D(net_2656), .CK(net_16725) );
CLKBUF_X2 inst_17179 ( .A(net_10166), .Z(net_17027) );
INV_X8 inst_5035 ( .ZN(net_6091), .A(net_3559) );
NAND2_X2 inst_4759 ( .ZN(net_5983), .A1(net_2008), .A2(net_1730) );
SDFFR_X2 inst_2392 ( .SE(net_2260), .Q(net_356), .D(net_356), .CK(net_10411), .RN(x6501), .SI(x2068) );
NAND2_X2 inst_4678 ( .A1(net_6114), .ZN(net_2580), .A2(net_2090) );
CLKBUF_X2 inst_9531 ( .A(net_9378), .Z(net_9379) );
NAND4_X2 inst_3667 ( .A4(net_6042), .A1(net_6041), .ZN(net_4598), .A2(net_4090), .A3(net_4089) );
CLKBUF_X2 inst_13513 ( .A(net_13360), .Z(net_13361) );
AOI22_X2 inst_7972 ( .B1(net_8195), .A1(net_7685), .B2(net_6099), .A2(net_4399), .ZN(net_4157) );
NAND2_X2 inst_4434 ( .A1(net_6871), .A2(net_5016), .ZN(net_4993) );
CLKBUF_X2 inst_14775 ( .A(net_14622), .Z(net_14623) );
CLKBUF_X2 inst_18841 ( .A(net_12449), .Z(net_18689) );
INV_X2 inst_6380 ( .ZN(net_1602), .A(net_1348) );
MUX2_X2 inst_4967 ( .A(net_7394), .S(net_2378), .Z(net_2356), .B(net_802) );
DFFR_X2 inst_7217 ( .QN(net_6410), .D(net_2337), .CK(net_18001), .RN(x6501) );
CLKBUF_X2 inst_14953 ( .A(net_14800), .Z(net_14801) );
DFF_X1 inst_6785 ( .Q(net_7534), .D(net_4585), .CK(net_11958) );
CLKBUF_X2 inst_10792 ( .A(net_10639), .Z(net_10640) );
SDFF_X2 inst_656 ( .Q(net_8428), .D(net_8428), .SI(net_3957), .SE(net_3934), .CK(net_13255) );
CLKBUF_X2 inst_10866 ( .A(net_10713), .Z(net_10714) );
CLKBUF_X2 inst_13993 ( .A(net_13840), .Z(net_13841) );
DFFS_X2 inst_6900 ( .QN(net_7160), .D(net_2326), .CK(net_15081), .SN(x6501) );
CLKBUF_X2 inst_9690 ( .A(net_9447), .Z(net_9538) );
XOR2_X2 inst_45 ( .A(net_6828), .B(net_1221), .Z(net_1036) );
CLKBUF_X2 inst_15351 ( .A(net_15198), .Z(net_15199) );
CLKBUF_X2 inst_9551 ( .A(net_9398), .Z(net_9399) );
CLKBUF_X2 inst_12500 ( .A(net_12347), .Z(net_12348) );
CLKBUF_X2 inst_15125 ( .A(net_9106), .Z(net_14973) );
SDFF_X2 inst_458 ( .SI(net_8461), .Q(net_8461), .SE(net_3983), .D(net_3944), .CK(net_12285) );
OAI21_X2 inst_3093 ( .B2(net_2861), .ZN(net_2860), .B1(net_1786), .A(net_1714) );
SDFF_X2 inst_1562 ( .Q(net_8027), .D(net_8027), .SI(net_2719), .SE(net_2545), .CK(net_16048) );
CLKBUF_X2 inst_9934 ( .A(net_9781), .Z(net_9782) );
NAND2_X2 inst_4148 ( .ZN(net_5369), .A1(net_5211), .A2(net_4998) );
CLKBUF_X2 inst_11814 ( .A(net_11114), .Z(net_11662) );
CLKBUF_X2 inst_17407 ( .A(net_9843), .Z(net_17255) );
INV_X4 inst_5539 ( .A(net_943), .ZN(net_865) );
AOI222_X1 inst_8644 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3924), .B1(net_3196), .C1(net_3194), .A1(x13815) );
SDFF_X2 inst_741 ( .Q(net_8782), .D(net_8782), .SI(net_3938), .SE(net_3879), .CK(net_12956) );
CLKBUF_X2 inst_18440 ( .A(net_18287), .Z(net_18288) );
CLKBUF_X2 inst_18063 ( .A(net_17910), .Z(net_17911) );
CLKBUF_X2 inst_9377 ( .A(net_9224), .Z(net_9225) );
CLKBUF_X2 inst_16976 ( .A(net_16823), .Z(net_16824) );
DFFR_X2 inst_7195 ( .QN(net_8956), .D(net_2421), .CK(net_15061), .RN(x6501) );
AOI222_X1 inst_8700 ( .B2(net_4889), .A2(net_4888), .C2(net_4803), .ZN(net_2937), .A1(net_2936), .B1(net_2935), .C1(net_858) );
CLKBUF_X2 inst_9338 ( .A(net_9130), .Z(net_9186) );
CLKBUF_X2 inst_10178 ( .A(net_9716), .Z(net_10026) );
CLKBUF_X2 inst_12964 ( .A(net_12811), .Z(net_12812) );
AOI22_X2 inst_8124 ( .B1(net_8014), .A1(net_7980), .B2(net_6102), .A2(net_6097), .ZN(net_4025) );
CLKBUF_X2 inst_17349 ( .A(net_17196), .Z(net_17197) );
OR2_X4 inst_2828 ( .ZN(net_3528), .A2(net_3527), .A1(net_3526) );
AOI22_X2 inst_7769 ( .B1(net_6996), .A1(net_6956), .A2(net_5443), .B2(net_5442), .ZN(net_5328) );
CLKBUF_X2 inst_13560 ( .A(net_9508), .Z(net_13408) );
NAND2_X2 inst_4745 ( .ZN(net_2589), .A2(net_1586), .A1(net_1462) );
NAND3_X4 inst_3877 ( .A3(net_7343), .ZN(net_6106), .A1(net_6094), .A2(net_718) );
CLKBUF_X2 inst_9859 ( .A(net_9706), .Z(net_9707) );
CLKBUF_X2 inst_16236 ( .A(net_16083), .Z(net_16084) );
CLKBUF_X2 inst_17300 ( .A(net_11948), .Z(net_17148) );
DFFR_X2 inst_7320 ( .QN(net_6466), .D(net_6463), .CK(net_15088), .RN(x6501) );
SDFF_X2 inst_1131 ( .D(net_7338), .SI(net_6580), .Q(net_6580), .SE(net_3070), .CK(net_9450) );
CLKBUF_X2 inst_14617 ( .A(net_14464), .Z(net_14465) );
SDFF_X2 inst_691 ( .Q(net_8886), .D(net_8886), .SI(net_3939), .SE(net_3936), .CK(net_12532) );
CLKBUF_X2 inst_14538 ( .A(net_14385), .Z(net_14386) );
CLKBUF_X2 inst_18523 ( .A(net_18370), .Z(net_18371) );
CLKBUF_X2 inst_11769 ( .A(net_10070), .Z(net_11617) );
INV_X2 inst_6402 ( .ZN(net_1592), .A(net_622) );
CLKBUF_X2 inst_12845 ( .A(net_12692), .Z(net_12693) );
SDFF_X2 inst_770 ( .Q(net_8814), .D(net_8814), .SI(net_3948), .SE(net_3879), .CK(net_13466) );
SDFF_X2 inst_565 ( .Q(net_8828), .D(net_8828), .SI(net_3966), .SE(net_3964), .CK(net_10015) );
CLKBUF_X2 inst_15912 ( .A(net_10545), .Z(net_15760) );
SDFF_X2 inst_622 ( .SI(net_8533), .Q(net_8533), .SE(net_3979), .D(net_3959), .CK(net_13194) );
SDFF_X2 inst_1971 ( .D(net_7282), .SI(net_6899), .Q(net_6899), .SE(net_6284), .CK(net_16165) );
DFFR_X1 inst_7418 ( .D(net_5581), .CK(net_13895), .RN(x6501), .Q(x641) );
CLKBUF_X2 inst_12342 ( .A(net_12189), .Z(net_12190) );
CLKBUF_X2 inst_14345 ( .A(net_14192), .Z(net_14193) );
CLKBUF_X2 inst_17772 ( .A(net_15094), .Z(net_17620) );
CLKBUF_X2 inst_17206 ( .A(net_17053), .Z(net_17054) );
CLKBUF_X2 inst_14531 ( .A(net_14378), .Z(net_14379) );
SDFF_X2 inst_409 ( .SI(net_8323), .Q(net_8323), .SE(net_3978), .D(net_3975), .CK(net_12555) );
CLKBUF_X2 inst_11679 ( .A(net_9549), .Z(net_11527) );
CLKBUF_X2 inst_12323 ( .A(net_10935), .Z(net_12171) );
CLKBUF_X2 inst_17181 ( .A(net_17028), .Z(net_17029) );
HA_X1 inst_6672 ( .A(net_7512), .CO(net_3263), .S(net_3197), .B(net_3007) );
INV_X4 inst_5813 ( .A(net_7496), .ZN(net_3056) );
CLKBUF_X2 inst_15611 ( .A(net_15458), .Z(net_15459) );
AOI22_X2 inst_8013 ( .B1(net_8166), .A1(net_7724), .B2(net_6101), .A2(net_6095), .ZN(net_4122) );
CLKBUF_X2 inst_12933 ( .A(net_12780), .Z(net_12781) );
NOR2_X2 inst_3506 ( .A1(net_3023), .ZN(net_1848), .A2(net_1671) );
CLKBUF_X2 inst_17478 ( .A(net_17325), .Z(net_17326) );
CLKBUF_X2 inst_9220 ( .A(net_9067), .Z(net_9068) );
CLKBUF_X2 inst_18880 ( .A(net_18727), .Z(net_18728) );
DFFR_X1 inst_7396 ( .D(net_5837), .CK(net_17172), .RN(x6501), .Q(x186) );
DFFR_X2 inst_7092 ( .QN(net_8292), .D(net_3551), .CK(net_11235), .RN(x6501) );
CLKBUF_X2 inst_11947 ( .A(net_11794), .Z(net_11795) );
CLKBUF_X2 inst_11389 ( .A(net_11236), .Z(net_11237) );
AOI22_X2 inst_7795 ( .A2(net_6187), .B2(net_5609), .ZN(net_4794), .B1(net_370), .A1(net_194) );
CLKBUF_X2 inst_15198 ( .A(net_15045), .Z(net_15046) );
SDFF_X2 inst_663 ( .Q(net_8410), .D(net_8410), .SI(net_3980), .SE(net_3934), .CK(net_10720) );
NOR4_X2 inst_3227 ( .ZN(net_3181), .A3(net_2309), .A4(net_2308), .A1(net_2244), .A2(net_1705) );
AOI21_X2 inst_8949 ( .A(net_5746), .ZN(net_5671), .B2(net_5451), .B1(net_4966) );
CLKBUF_X2 inst_16493 ( .A(net_16340), .Z(net_16341) );
NAND2_X2 inst_4224 ( .A1(net_7016), .A2(net_5249), .ZN(net_5236) );
DFFR_X2 inst_7279 ( .QN(net_6391), .D(net_1848), .CK(net_15664), .RN(x6501) );
SDFFR_X2 inst_2290 ( .SI(net_2475), .SE(net_2426), .Q(net_434), .D(net_434), .CK(net_16422), .RN(x6501) );
CLKBUF_X2 inst_17463 ( .A(net_15738), .Z(net_17311) );
CLKBUF_X2 inst_11913 ( .A(net_11760), .Z(net_11761) );
INV_X4 inst_5070 ( .ZN(net_5858), .A(net_5812) );
INV_X4 inst_5797 ( .A(net_6345), .ZN(net_744) );
CLKBUF_X2 inst_14640 ( .A(net_14487), .Z(net_14488) );
SDFFR_X2 inst_2621 ( .Q(net_7390), .D(net_7390), .SE(net_1136), .CK(net_18311), .RN(x6501), .SI(x4538) );
CLKBUF_X2 inst_15743 ( .A(net_15590), .Z(net_15591) );
AND2_X2 inst_9159 ( .ZN(net_2811), .A1(net_2810), .A2(net_2809) );
CLKBUF_X2 inst_10815 ( .A(net_10169), .Z(net_10663) );
CLKBUF_X2 inst_14454 ( .A(net_14301), .Z(net_14302) );
CLKBUF_X2 inst_18559 ( .A(net_14187), .Z(net_18407) );
CLKBUF_X2 inst_16598 ( .A(net_16445), .Z(net_16446) );
CLKBUF_X2 inst_11928 ( .A(net_9603), .Z(net_11776) );
CLKBUF_X2 inst_9358 ( .A(net_9205), .Z(net_9206) );
SDFF_X2 inst_1647 ( .SI(net_7726), .Q(net_7726), .D(net_2712), .SE(net_2559), .CK(net_13770) );
NOR3_X2 inst_3263 ( .ZN(net_3021), .A1(net_2975), .A3(net_877), .A2(net_506) );
CLKBUF_X2 inst_12114 ( .A(net_11961), .Z(net_11962) );
SDFF_X2 inst_1376 ( .SI(net_7276), .Q(net_7133), .D(net_7133), .SE(net_6279), .CK(net_17401) );
OR2_X2 inst_2882 ( .A2(net_9008), .A1(net_6118), .ZN(net_2262) );
CLKBUF_X2 inst_10507 ( .A(net_9365), .Z(net_10355) );
CLKBUF_X2 inst_12605 ( .A(net_12452), .Z(net_12453) );
CLKBUF_X2 inst_18325 ( .A(net_18172), .Z(net_18173) );
AOI22_X2 inst_8182 ( .B1(net_8753), .A1(net_8383), .A2(net_3867), .B2(net_3866), .ZN(net_3850) );
CLKBUF_X2 inst_11483 ( .A(net_11330), .Z(net_11331) );
CLKBUF_X2 inst_10654 ( .A(net_10501), .Z(net_10502) );
INV_X2 inst_6188 ( .ZN(net_5793), .A(net_5759) );
CLKBUF_X2 inst_10742 ( .A(net_10148), .Z(net_10590) );
SDFF_X2 inst_1659 ( .SI(net_7749), .Q(net_7749), .D(net_2706), .SE(net_2560), .CK(net_18850) );
CLKBUF_X2 inst_17331 ( .A(net_17178), .Z(net_17179) );
AOI22_X2 inst_8184 ( .B1(net_8790), .A1(net_8531), .A2(net_3861), .B2(net_3860), .ZN(net_3848) );
INV_X4 inst_5702 ( .A(net_7237), .ZN(net_1952) );
SDFF_X2 inst_398 ( .SI(net_8310), .Q(net_8310), .SE(net_3978), .D(net_3966), .CK(net_10943) );
SDFF_X2 inst_436 ( .Q(net_8764), .D(net_8764), .SE(net_3982), .SI(net_3942), .CK(net_12640) );
CLKBUF_X2 inst_11766 ( .A(net_11613), .Z(net_11614) );
CLKBUF_X2 inst_13265 ( .A(net_13112), .Z(net_13113) );
INV_X2 inst_6529 ( .A(net_7493), .ZN(net_523) );
CLKBUF_X2 inst_9852 ( .A(net_9511), .Z(net_9700) );
NAND4_X2 inst_3705 ( .ZN(net_4432), .A4(net_4336), .A1(net_3733), .A2(net_3732), .A3(net_3731) );
CLKBUF_X2 inst_19077 ( .A(net_18924), .Z(net_18925) );
CLKBUF_X2 inst_17990 ( .A(net_17837), .Z(net_17838) );
DFF_X1 inst_6746 ( .QN(net_6790), .D(net_5623), .CK(net_11580) );
SDFFR_X2 inst_2231 ( .Q(net_7464), .D(net_7464), .SE(net_2863), .CK(net_12167), .SI(x13482), .RN(x6501) );
XNOR2_X2 inst_144 ( .ZN(net_2289), .B(net_2017), .A(net_1828) );
CLKBUF_X2 inst_18891 ( .A(net_18738), .Z(net_18739) );
CLKBUF_X2 inst_9750 ( .A(net_9597), .Z(net_9598) );
CLKBUF_X2 inst_10565 ( .A(net_10412), .Z(net_10413) );
CLKBUF_X2 inst_13660 ( .A(net_13507), .Z(net_13508) );
CLKBUF_X2 inst_18230 ( .A(net_18077), .Z(net_18078) );
DFFS_X1 inst_6912 ( .D(net_5736), .CK(net_13813), .SN(x6501), .Q(x0) );
CLKBUF_X2 inst_17524 ( .A(net_17371), .Z(net_17372) );
NAND2_X2 inst_4857 ( .A1(net_8214), .ZN(net_1152), .A2(net_742) );
CLKBUF_X2 inst_9763 ( .A(net_9610), .Z(net_9611) );
CLKBUF_X2 inst_16892 ( .A(net_16739), .Z(net_16740) );
INV_X4 inst_5555 ( .A(net_1459), .ZN(net_634) );
CLKBUF_X2 inst_10026 ( .A(net_9495), .Z(net_9874) );
NAND2_X2 inst_4447 ( .A1(net_6847), .A2(net_5016), .ZN(net_4980) );
INV_X2 inst_6194 ( .A(net_6789), .ZN(net_5732) );
AOI22_X2 inst_8493 ( .B1(net_6745), .A1(net_6712), .B2(net_6202), .A2(net_3520), .ZN(net_3447) );
CLKBUF_X2 inst_15694 ( .A(net_15541), .Z(net_15542) );
CLKBUF_X2 inst_17818 ( .A(net_14625), .Z(net_17666) );
INV_X2 inst_6329 ( .A(net_3296), .ZN(net_3174) );
CLKBUF_X2 inst_12470 ( .A(net_12317), .Z(net_12318) );
CLKBUF_X2 inst_16065 ( .A(net_15912), .Z(net_15913) );
CLKBUF_X2 inst_15878 ( .A(net_15725), .Z(net_15726) );
CLKBUF_X2 inst_14937 ( .A(net_11093), .Z(net_14785) );
SDFF_X2 inst_1360 ( .Q(net_8202), .D(net_8202), .SI(net_2712), .SE(net_2561), .CK(net_17148) );
CLKBUF_X2 inst_15871 ( .A(net_15718), .Z(net_15719) );
CLKBUF_X2 inst_16578 ( .A(net_15065), .Z(net_16426) );
SDFF_X2 inst_466 ( .SI(net_8471), .Q(net_8471), .SE(net_3983), .D(net_3975), .CK(net_12552) );
NAND3_X2 inst_3981 ( .A2(net_2530), .A1(net_2250), .ZN(net_2216), .A3(net_1899) );
CLKBUF_X2 inst_18237 ( .A(net_18084), .Z(net_18085) );
INV_X4 inst_5205 ( .A(net_5718), .ZN(net_2395) );
CLKBUF_X2 inst_14742 ( .A(net_10930), .Z(net_14590) );
CLKBUF_X2 inst_10073 ( .A(net_9920), .Z(net_9921) );
OAI21_X2 inst_3038 ( .B2(net_8241), .B1(net_4928), .ZN(net_4840), .A(net_3335) );
CLKBUF_X2 inst_14154 ( .A(net_13557), .Z(net_14002) );
DFFR_X1 inst_7542 ( .D(net_2698), .Q(net_290), .CK(net_9667), .RN(x6501) );
CLKBUF_X2 inst_16863 ( .A(net_16710), .Z(net_16711) );
NAND3_X4 inst_3864 ( .A3(net_6259), .A1(net_6193), .ZN(net_4904), .A2(net_4901) );
CLKBUF_X2 inst_15482 ( .A(net_15329), .Z(net_15330) );
CLKBUF_X2 inst_12735 ( .A(net_12582), .Z(net_12583) );
CLKBUF_X2 inst_15596 ( .A(net_15443), .Z(net_15444) );
DFFR_X1 inst_7406 ( .D(net_5706), .CK(net_14043), .RN(x6501), .Q(x378) );
CLKBUF_X2 inst_9757 ( .A(net_9604), .Z(net_9605) );
CLKBUF_X2 inst_18566 ( .A(net_18413), .Z(net_18414) );
DFFR_X2 inst_7283 ( .QN(net_7523), .D(net_1721), .CK(net_16289), .RN(x6501) );
INV_X4 inst_5214 ( .ZN(net_2945), .A(net_2338) );
CLKBUF_X2 inst_15170 ( .A(net_15017), .Z(net_15018) );
CLKBUF_X2 inst_13331 ( .A(net_13178), .Z(net_13179) );
NAND2_X2 inst_4794 ( .A1(net_2255), .ZN(net_1482), .A2(net_1132) );
CLKBUF_X2 inst_13838 ( .A(net_13685), .Z(net_13686) );
CLKBUF_X2 inst_10804 ( .A(net_10651), .Z(net_10652) );
CLKBUF_X2 inst_13688 ( .A(net_13535), .Z(net_13536) );
NAND4_X2 inst_3829 ( .A4(net_6258), .ZN(net_2963), .A3(net_1282), .A1(net_1091), .A2(net_265) );
AOI22_X2 inst_7883 ( .B1(net_7196), .A2(net_6447), .B2(net_5655), .A1(net_5654), .ZN(net_4548) );
CLKBUF_X2 inst_14465 ( .A(net_12740), .Z(net_14313) );
CLKBUF_X2 inst_17755 ( .A(net_17602), .Z(net_17603) );
AOI211_X2 inst_9012 ( .C2(net_6187), .ZN(net_4935), .A(net_4834), .B(net_4658), .C1(net_187) );
CLKBUF_X2 inst_13414 ( .A(net_13261), .Z(net_13262) );
CLKBUF_X2 inst_14621 ( .A(net_14468), .Z(net_14469) );
CLKBUF_X2 inst_10325 ( .A(net_10172), .Z(net_10173) );
CLKBUF_X2 inst_10971 ( .A(net_10818), .Z(net_10819) );
CLKBUF_X2 inst_13918 ( .A(net_13765), .Z(net_13766) );
CLKBUF_X2 inst_15791 ( .A(net_14910), .Z(net_15639) );
CLKBUF_X2 inst_17811 ( .A(net_17658), .Z(net_17659) );
AOI22_X2 inst_8161 ( .B1(net_8852), .A1(net_8297), .B2(net_6252), .A2(net_4345), .ZN(net_3873) );
SDFFR_X2 inst_2168 ( .QN(net_7592), .D(net_3951), .SE(net_3144), .SI(net_3134), .CK(net_10388), .RN(x6501) );
DFFR_X2 inst_7241 ( .QN(net_5957), .D(net_2057), .CK(net_15058), .RN(x6501) );
CLKBUF_X2 inst_15060 ( .A(net_14907), .Z(net_14908) );
CLKBUF_X2 inst_18889 ( .A(net_18736), .Z(net_18737) );
NAND2_X2 inst_4322 ( .A1(net_7059), .A2(net_5162), .ZN(net_5135) );
SDFF_X2 inst_1078 ( .D(net_7329), .SI(net_6505), .Q(net_6505), .SE(net_3071), .CK(net_9513) );
INV_X2 inst_6497 ( .ZN(net_3018), .A(x13291) );
NOR2_X2 inst_3557 ( .ZN(net_1503), .A1(net_825), .A2(net_602) );
SDFF_X2 inst_1039 ( .SI(net_7337), .Q(net_6711), .D(net_6711), .SE(net_3125), .CK(net_9484) );
SDFF_X2 inst_1992 ( .SI(net_7912), .Q(net_7912), .D(net_2709), .SE(net_2461), .CK(net_15810) );
CLKBUF_X2 inst_16679 ( .A(net_12085), .Z(net_16527) );
INV_X4 inst_5449 ( .A(net_1633), .ZN(net_1148) );
NAND2_X4 inst_4048 ( .A1(net_6106), .A2(net_2185), .ZN(net_2170) );
DFFR_X1 inst_7549 ( .Q(net_7641), .D(net_577), .CK(net_15706), .RN(x6501) );
NAND3_X2 inst_4003 ( .A1(net_7401), .A3(net_1504), .ZN(net_1432), .A2(net_670) );
DFFS_X2 inst_6868 ( .QN(net_6807), .D(net_4623), .CK(net_11805), .SN(x6501) );
INV_X8 inst_5033 ( .ZN(net_2299), .A(net_2187) );
AOI22_X2 inst_8306 ( .A1(net_8622), .B1(net_8437), .A2(net_3864), .B2(net_3863), .ZN(net_3739) );
CLKBUF_X2 inst_15512 ( .A(net_15359), .Z(net_15360) );
CLKBUF_X2 inst_13966 ( .A(net_13160), .Z(net_13814) );
AOI221_X2 inst_8846 ( .B1(net_8567), .C1(net_8456), .C2(net_6263), .B2(net_6262), .ZN(net_6243), .A(net_4265) );
INV_X4 inst_5363 ( .ZN(net_1344), .A(net_757) );
CLKBUF_X2 inst_17128 ( .A(net_11952), .Z(net_16976) );
NOR2_X2 inst_3542 ( .ZN(net_2247), .A2(net_1669), .A1(net_1475) );
CLKBUF_X2 inst_15529 ( .A(net_15376), .Z(net_15377) );
CLKBUF_X2 inst_16547 ( .A(net_16394), .Z(net_16395) );
INV_X2 inst_6300 ( .ZN(net_4023), .A(net_3907) );
XNOR2_X2 inst_115 ( .B(net_7513), .ZN(net_6214), .A(net_3264) );
NAND2_X2 inst_4691 ( .ZN(net_4821), .A1(net_4320), .A2(net_2066) );
NAND4_X2 inst_3726 ( .ZN(net_4304), .A2(net_4160), .A1(net_4159), .A3(net_4158), .A4(net_4157) );
OAI21_X2 inst_3045 ( .B2(net_8227), .B1(net_4928), .ZN(net_4776), .A(net_2970) );
CLKBUF_X2 inst_9801 ( .A(net_9648), .Z(net_9649) );
CLKBUF_X2 inst_12741 ( .A(net_10468), .Z(net_12589) );
CLKBUF_X2 inst_18877 ( .A(net_18043), .Z(net_18725) );
INV_X4 inst_6113 ( .A(net_7574), .ZN(net_485) );
SDFF_X2 inst_1263 ( .Q(net_8108), .D(net_8108), .SE(net_2707), .SI(net_2704), .CK(net_17032) );
CLKBUF_X2 inst_16699 ( .A(net_16546), .Z(net_16547) );
AOI22_X2 inst_8047 ( .B1(net_7933), .A1(net_7831), .B2(net_6103), .A2(net_4398), .ZN(net_4093) );
NOR2_X4 inst_3330 ( .ZN(net_3369), .A2(net_3180), .A1(net_3119) );
CLKBUF_X2 inst_10225 ( .A(net_10072), .Z(net_10073) );
DFFR_X1 inst_7374 ( .QN(net_5944), .D(net_5887), .CK(net_9407), .RN(x6501) );
SDFF_X2 inst_1445 ( .SI(net_7265), .Q(net_7082), .D(net_7082), .SE(net_6278), .CK(net_17079) );
CLKBUF_X2 inst_11907 ( .A(net_11754), .Z(net_11755) );
CLKBUF_X2 inst_16728 ( .A(net_16575), .Z(net_16576) );
NAND3_X2 inst_3990 ( .A2(net_9047), .ZN(net_3950), .A1(net_1593), .A3(net_1592) );
CLKBUF_X2 inst_17500 ( .A(net_15852), .Z(net_17348) );
AOI21_X2 inst_8976 ( .A(net_2222), .ZN(net_2191), .B2(net_2187), .B1(net_919) );
CLKBUF_X2 inst_18318 ( .A(net_18165), .Z(net_18166) );
CLKBUF_X2 inst_13156 ( .A(net_13003), .Z(net_13004) );
INV_X4 inst_5982 ( .A(net_6381), .ZN(net_1492) );
CLKBUF_X2 inst_12115 ( .A(net_11962), .Z(net_11963) );
AOI22_X2 inst_7931 ( .B1(net_8054), .A1(net_7850), .B2(net_6107), .ZN(net_5998), .A2(net_4400) );
CLKBUF_X2 inst_15945 ( .A(net_9341), .Z(net_15793) );
CLKBUF_X2 inst_16744 ( .A(net_16591), .Z(net_16592) );
AOI22_X2 inst_7932 ( .A1(net_7952), .B1(net_7782), .A2(net_6092), .B2(net_6091), .ZN(net_4193) );
SDFF_X2 inst_1512 ( .SI(net_7873), .Q(net_7873), .D(net_2703), .SE(net_2558), .CK(net_14014) );
CLKBUF_X2 inst_10366 ( .A(net_10213), .Z(net_10214) );
INV_X4 inst_5160 ( .ZN(net_5835), .A(net_3059) );
AOI221_X4 inst_8733 ( .B1(net_8739), .C1(net_8517), .B2(net_4350), .C2(net_4349), .ZN(net_4333), .A(net_4239) );
CLKBUF_X2 inst_13209 ( .A(net_9349), .Z(net_13057) );
CLKBUF_X2 inst_14395 ( .A(net_14242), .Z(net_14243) );
CLKBUF_X2 inst_18791 ( .A(net_18638), .Z(net_18639) );
CLKBUF_X2 inst_10727 ( .A(net_9451), .Z(net_10575) );
CLKBUF_X2 inst_16017 ( .A(net_13617), .Z(net_15865) );
CLKBUF_X2 inst_14822 ( .A(net_14669), .Z(net_14670) );
SDFFR_X2 inst_2299 ( .D(net_2968), .SE(net_2313), .SI(net_410), .Q(net_410), .CK(net_13957), .RN(x6501) );
CLKBUF_X2 inst_11691 ( .A(net_11538), .Z(net_11539) );
CLKBUF_X2 inst_12441 ( .A(net_12288), .Z(net_12289) );
CLKBUF_X2 inst_19184 ( .A(net_19031), .Z(net_19032) );
DFFR_X1 inst_7504 ( .Q(net_7222), .D(net_2074), .CK(net_15217), .RN(x6501) );
INV_X4 inst_5292 ( .ZN(net_1606), .A(net_1605) );
CLKBUF_X2 inst_16829 ( .A(net_9677), .Z(net_16677) );
DFFR_X1 inst_7578 ( .D(x192486), .Q(net_384), .CK(net_18730), .RN(x6501) );
AOI22_X2 inst_8166 ( .A1(net_8593), .B1(net_8408), .ZN(net_3870), .A2(net_3864), .B2(net_3863) );
CLKBUF_X2 inst_12366 ( .A(net_11705), .Z(net_12214) );
CLKBUF_X2 inst_14963 ( .A(net_14810), .Z(net_14811) );
SDFF_X2 inst_1642 ( .SI(net_7716), .Q(net_7716), .D(net_2574), .SE(net_2559), .CK(net_16037) );
CLKBUF_X2 inst_12703 ( .A(net_12550), .Z(net_12551) );
CLKBUF_X2 inst_13434 ( .A(net_13281), .Z(net_13282) );
XNOR2_X2 inst_199 ( .ZN(net_1545), .B(net_1195), .A(net_1190) );
CLKBUF_X2 inst_12540 ( .A(net_12387), .Z(net_12388) );
CLKBUF_X2 inst_13259 ( .A(net_13106), .Z(net_13107) );
DFF_X1 inst_6764 ( .Q(net_7544), .D(net_4608), .CK(net_9728) );
DFFR_X2 inst_6976 ( .QN(net_5975), .D(net_5901), .CK(net_11559), .RN(x6501) );
CLKBUF_X2 inst_13313 ( .A(net_13160), .Z(net_13161) );
NAND2_X2 inst_4875 ( .A2(net_3334), .ZN(net_1153), .A1(net_477) );
CLKBUF_X2 inst_14274 ( .A(net_14121), .Z(net_14122) );
CLKBUF_X2 inst_16956 ( .A(net_16803), .Z(net_16804) );
CLKBUF_X2 inst_18163 ( .A(net_18010), .Z(net_18011) );
CLKBUF_X2 inst_14252 ( .A(net_11203), .Z(net_14100) );
CLKBUF_X2 inst_15412 ( .A(net_15259), .Z(net_15260) );
NAND2_X2 inst_4114 ( .ZN(net_5415), .A2(net_5234), .A1(net_5141) );
SDFF_X2 inst_540 ( .Q(net_8682), .D(net_8682), .SI(net_3973), .SE(net_3935), .CK(net_12342) );
SDFFR_X2 inst_2356 ( .SE(net_2313), .D(net_719), .SI(net_463), .Q(net_463), .CK(net_16731), .RN(x6501) );
SDFF_X2 inst_998 ( .D(net_7338), .SI(net_6646), .Q(net_6646), .SE(net_3123), .CK(net_9496) );
AOI22_X2 inst_7989 ( .B1(net_8096), .A1(net_7756), .B2(net_6108), .A2(net_6096), .ZN(net_4143) );
INV_X4 inst_6044 ( .A(net_7485), .ZN(net_2290) );
INV_X4 inst_5952 ( .A(net_7609), .ZN(net_2752) );
OAI211_X2 inst_3209 ( .ZN(net_2174), .B(net_1905), .C2(net_1904), .A(net_1723), .C1(net_1722) );
CLKBUF_X2 inst_13989 ( .A(net_13836), .Z(net_13837) );
CLKBUF_X2 inst_9730 ( .A(net_9577), .Z(net_9578) );
CLKBUF_X2 inst_12298 ( .A(net_12145), .Z(net_12146) );
CLKBUF_X2 inst_14042 ( .A(net_12520), .Z(net_13890) );
CLKBUF_X2 inst_9792 ( .A(net_9639), .Z(net_9640) );
CLKBUF_X2 inst_9242 ( .A(net_9089), .Z(net_9090) );
CLKBUF_X2 inst_10205 ( .A(net_10052), .Z(net_10053) );
CLKBUF_X2 inst_11442 ( .A(net_11289), .Z(net_11290) );
INV_X4 inst_5090 ( .ZN(net_5707), .A(net_5684) );
DFF_X1 inst_6720 ( .Q(net_6766), .D(net_5649), .CK(net_9273) );
XNOR2_X2 inst_192 ( .A(net_7659), .ZN(net_1554), .B(net_1553) );
CLKBUF_X2 inst_14400 ( .A(net_14247), .Z(net_14248) );
SDFFR_X1 inst_2715 ( .SI(net_8891), .Q(net_7634), .D(net_7634), .SE(net_3901), .CK(net_13516), .RN(x6501) );
NAND2_X2 inst_4242 ( .A1(net_7024), .A2(net_5249), .ZN(net_5218) );
CLKBUF_X2 inst_13059 ( .A(net_12906), .Z(net_12907) );
NAND2_X2 inst_4126 ( .ZN(net_5399), .A2(net_5226), .A1(net_5129) );
DFFR_X1 inst_7434 ( .QN(net_8914), .D(net_4852), .CK(net_13981), .RN(x6501) );
NAND2_X2 inst_4178 ( .ZN(net_5326), .A1(net_5191), .A2(net_4988) );
NOR2_X2 inst_3547 ( .A1(net_1450), .ZN(net_1445), .A2(net_1064) );
AOI221_X2 inst_8741 ( .B2(net_8246), .ZN(net_5690), .A(net_5537), .B1(net_5268), .C2(net_5267), .C1(net_183) );
CLKBUF_X2 inst_12720 ( .A(net_12567), .Z(net_12568) );
INV_X2 inst_6558 ( .A(net_7568), .ZN(net_3110) );
CLKBUF_X2 inst_18901 ( .A(net_18748), .Z(net_18749) );
CLKBUF_X2 inst_9739 ( .A(net_9586), .Z(net_9587) );
DFFR_X2 inst_7234 ( .QN(net_6836), .D(net_2193), .CK(net_18724), .RN(x6501) );
SDFF_X2 inst_486 ( .SI(net_8609), .Q(net_8609), .SE(net_3984), .D(net_3944), .CK(net_10847) );
CLKBUF_X2 inst_12977 ( .A(net_12824), .Z(net_12825) );
CLKBUF_X2 inst_15117 ( .A(net_12104), .Z(net_14965) );
CLKBUF_X2 inst_13365 ( .A(net_9910), .Z(net_13213) );
SDFF_X2 inst_1240 ( .Q(net_7964), .D(net_7964), .SE(net_2755), .SI(net_2712), .CK(net_13799) );
INV_X4 inst_5445 ( .ZN(net_1082), .A(net_813) );
INV_X2 inst_6597 ( .ZN(net_6132), .A(net_6129) );
CLKBUF_X2 inst_18740 ( .A(net_18587), .Z(net_18588) );
CLKBUF_X2 inst_15941 ( .A(net_15788), .Z(net_15789) );
AND2_X2 inst_9186 ( .A2(net_2250), .ZN(net_2091), .A1(net_1900) );
SDFF_X2 inst_1521 ( .Q(net_7892), .D(net_7892), .SI(net_2590), .SE(net_2543), .CK(net_15598) );
INV_X2 inst_6620 ( .ZN(net_6256), .A(net_6255) );
CLKBUF_X2 inst_13692 ( .A(net_10877), .Z(net_13540) );
CLKBUF_X2 inst_9679 ( .A(net_9526), .Z(net_9527) );
CLKBUF_X2 inst_12976 ( .A(net_12823), .Z(net_12824) );
NAND2_X2 inst_4845 ( .ZN(net_1413), .A1(net_908), .A2(net_907) );
SDFF_X2 inst_1306 ( .Q(net_7818), .D(net_7818), .SE(net_2730), .SI(net_2574), .CK(net_17721) );
SDFFR_X2 inst_2563 ( .SI(net_7262), .Q(net_7262), .D(net_2127), .SE(net_1379), .CK(net_15031), .RN(x6501) );
CLKBUF_X2 inst_10766 ( .A(net_10613), .Z(net_10614) );
CLKBUF_X2 inst_11208 ( .A(net_10073), .Z(net_11056) );
CLKBUF_X2 inst_18007 ( .A(net_17854), .Z(net_17855) );
CLKBUF_X2 inst_9931 ( .A(net_9656), .Z(net_9779) );
CLKBUF_X2 inst_15640 ( .A(net_15487), .Z(net_15488) );
SDFF_X2 inst_1407 ( .SI(net_7275), .Q(net_7052), .D(net_7052), .SE(net_6280), .CK(net_17392) );
CLKBUF_X2 inst_12916 ( .A(net_12763), .Z(net_12764) );
AOI22_X2 inst_8096 ( .B1(net_8109), .A1(net_7769), .B2(net_6108), .A2(net_6096), .ZN(net_4051) );
CLKBUF_X2 inst_13128 ( .A(net_12975), .Z(net_12976) );
CLKBUF_X2 inst_13803 ( .A(net_11373), .Z(net_13651) );
DFFR_X2 inst_7018 ( .QN(net_9014), .D(net_5748), .CK(net_11171), .RN(x6501) );
CLKBUF_X2 inst_16176 ( .A(net_12806), .Z(net_16024) );
AND2_X4 inst_9132 ( .ZN(net_1401), .A2(net_815), .A1(net_171) );
INV_X4 inst_6052 ( .A(net_8895), .ZN(net_3187) );
CLKBUF_X2 inst_11526 ( .A(net_9644), .Z(net_11374) );
CLKBUF_X2 inst_17862 ( .A(net_17709), .Z(net_17710) );
DFFS_X1 inst_6965 ( .D(net_6829), .Q(net_6802), .CK(net_9632), .SN(x6501) );
CLKBUF_X2 inst_11051 ( .A(net_10898), .Z(net_10899) );
CLKBUF_X2 inst_9687 ( .A(net_9082), .Z(net_9535) );
CLKBUF_X2 inst_10217 ( .A(net_10064), .Z(net_10065) );
INV_X4 inst_5099 ( .ZN(net_5694), .A(net_5665) );
CLKBUF_X2 inst_11116 ( .A(net_10963), .Z(net_10964) );
INV_X4 inst_6134 ( .A(net_7580), .ZN(net_479) );
SDFF_X2 inst_584 ( .Q(net_8851), .D(net_8851), .SE(net_3964), .SI(net_3948), .CK(net_13415) );
CLKBUF_X2 inst_9561 ( .A(net_9106), .Z(net_9409) );
SDFF_X2 inst_470 ( .SI(net_8475), .Q(net_8475), .SE(net_3983), .D(net_3940), .CK(net_10282) );
AOI222_X1 inst_8668 ( .B1(net_7668), .A2(net_3599), .B2(net_3598), .C2(net_3597), .ZN(net_3590), .C1(net_1549), .A1(net_1182) );
CLKBUF_X2 inst_15566 ( .A(net_15413), .Z(net_15414) );
CLKBUF_X2 inst_12917 ( .A(net_12764), .Z(net_12765) );
AOI22_X2 inst_8138 ( .B1(net_8016), .A1(net_7982), .B2(net_6102), .A2(net_6097), .ZN(net_4012) );
NAND2_X2 inst_4490 ( .A1(net_7199), .A2(net_5655), .ZN(net_4482) );
SDFF_X2 inst_1752 ( .Q(net_8133), .D(net_8133), .SI(net_2713), .SE(net_2541), .CK(net_14391) );
CLKBUF_X2 inst_18221 ( .A(net_18068), .Z(net_18069) );
CLKBUF_X2 inst_16394 ( .A(net_16241), .Z(net_16242) );
DFF_X1 inst_6816 ( .QN(net_8231), .D(net_4450), .CK(net_14460) );
NAND2_X2 inst_4333 ( .A1(net_7102), .A2(net_5164), .ZN(net_5124) );
SDFF_X2 inst_1063 ( .D(net_7326), .SI(net_6634), .Q(net_6634), .SE(net_3123), .CK(net_11290) );
SDFFR_X1 inst_2700 ( .SI(net_7532), .SE(net_5043), .CK(net_11938), .RN(x6501), .Q(x4154), .D(x4154) );
NOR3_X2 inst_3252 ( .ZN(net_5737), .A2(net_5714), .A3(net_5712), .A1(net_5679) );
CLKBUF_X2 inst_13542 ( .A(net_13389), .Z(net_13390) );
NAND2_X2 inst_4565 ( .A1(net_6460), .A2(net_3294), .ZN(net_3121) );
NAND2_X2 inst_4755 ( .ZN(net_4510), .A1(net_2981), .A2(net_1733) );
CLKBUF_X2 inst_19100 ( .A(net_18947), .Z(net_18948) );
INV_X4 inst_5276 ( .A(net_2389), .ZN(net_1932) );
CLKBUF_X2 inst_18203 ( .A(net_18050), .Z(net_18051) );
CLKBUF_X2 inst_17375 ( .A(net_17222), .Z(net_17223) );
SDFF_X2 inst_1167 ( .D(net_7313), .SI(net_6489), .Q(net_6489), .SE(net_3071), .CK(net_11992) );
CLKBUF_X2 inst_9452 ( .A(net_9299), .Z(net_9300) );
DFFS_X2 inst_6879 ( .QN(net_6461), .D(net_3349), .CK(net_17922), .SN(x6501) );
CLKBUF_X2 inst_17931 ( .A(net_17778), .Z(net_17779) );
AOI221_X2 inst_8767 ( .C2(net_6131), .B2(net_5655), .ZN(net_5455), .A(net_4940), .B1(net_2955), .C1(net_1383) );
CLKBUF_X2 inst_14595 ( .A(net_14442), .Z(net_14443) );
SDFF_X2 inst_1303 ( .Q(net_8096), .D(net_8096), .SE(net_2707), .SI(net_2590), .CK(net_16006) );
SDFF_X2 inst_1623 ( .Q(net_8166), .D(net_8166), .SI(net_2718), .SE(net_2538), .CK(net_18777) );
NAND2_X2 inst_4088 ( .ZN(net_5581), .A2(net_5024), .A1(net_4958) );
CLKBUF_X2 inst_12788 ( .A(net_12635), .Z(net_12636) );
INV_X4 inst_6163 ( .A(net_6272), .ZN(net_6269) );
MUX2_X2 inst_4922 ( .S(net_6272), .A(net_6142), .Z(net_4618), .B(net_4617) );
AOI22_X2 inst_8369 ( .A1(net_8596), .B1(net_8411), .A2(net_3864), .B2(net_3863), .ZN(net_3679) );
NOR2_X2 inst_3452 ( .A1(net_3023), .ZN(net_2934), .A2(net_2825) );
CLKBUF_X2 inst_10183 ( .A(net_10030), .Z(net_10031) );
CLKBUF_X2 inst_17708 ( .A(net_10067), .Z(net_17556) );
SDFF_X2 inst_1516 ( .Q(net_7874), .D(net_7874), .SI(net_2721), .SE(net_2543), .CK(net_15843) );
CLKBUF_X2 inst_19047 ( .A(net_18894), .Z(net_18895) );
CLKBUF_X2 inst_14695 ( .A(net_10893), .Z(net_14543) );
SDFF_X2 inst_386 ( .Q(net_8822), .D(net_8822), .SI(net_3981), .SE(net_3964), .CK(net_10744) );
AOI22_X2 inst_8497 ( .B1(net_6746), .A1(net_6713), .B2(net_6202), .A2(net_3520), .ZN(net_3443) );
CLKBUF_X2 inst_12372 ( .A(net_10930), .Z(net_12220) );
CLKBUF_X2 inst_15110 ( .A(net_14957), .Z(net_14958) );
DFFR_X2 inst_7255 ( .QN(net_7234), .D(net_1982), .CK(net_17559), .RN(x6501) );
CLKBUF_X2 inst_10543 ( .A(net_10390), .Z(net_10391) );
CLKBUF_X2 inst_16914 ( .A(net_16761), .Z(net_16762) );
CLKBUF_X2 inst_9863 ( .A(net_9710), .Z(net_9711) );
CLKBUF_X2 inst_18780 ( .A(net_18627), .Z(net_18628) );
AOI22_X2 inst_8089 ( .B1(net_8108), .A1(net_7768), .B2(net_6108), .A2(net_6096), .ZN(net_4057) );
AOI22_X2 inst_7826 ( .A2(net_6430), .B2(net_5657), .A1(net_5654), .ZN(net_4696), .B1(net_2696) );
CLKBUF_X2 inst_11040 ( .A(net_10887), .Z(net_10888) );
CLKBUF_X2 inst_16220 ( .A(net_14931), .Z(net_16068) );
INV_X4 inst_5225 ( .A(net_2453), .ZN(net_2338) );
CLKBUF_X2 inst_16620 ( .A(net_16467), .Z(net_16468) );
INV_X4 inst_5320 ( .ZN(net_1662), .A(net_1301) );
SDFFR_X1 inst_2778 ( .Q(net_7292), .SI(net_1953), .D(net_1330), .SE(net_1327), .CK(net_15370), .RN(x6501) );
CLKBUF_X2 inst_9826 ( .A(net_9673), .Z(net_9674) );
CLKBUF_X2 inst_10173 ( .A(net_10020), .Z(net_10021) );
CLKBUF_X2 inst_11883 ( .A(net_11730), .Z(net_11731) );
INV_X4 inst_5223 ( .A(net_2453), .ZN(net_2281) );
INV_X4 inst_5468 ( .ZN(net_1323), .A(net_753) );
CLKBUF_X2 inst_19072 ( .A(net_18919), .Z(net_18920) );
CLKBUF_X2 inst_17265 ( .A(net_17112), .Z(net_17113) );
CLKBUF_X2 inst_9599 ( .A(net_9446), .Z(net_9447) );
AOI221_X4 inst_8716 ( .C1(net_7917), .B1(net_7815), .C2(net_6103), .ZN(net_6053), .B2(net_4398), .A(net_4277) );
CLKBUF_X2 inst_10060 ( .A(net_9907), .Z(net_9908) );
CLKBUF_X2 inst_11064 ( .A(net_10911), .Z(net_10912) );
SDFF_X2 inst_811 ( .SI(net_8501), .Q(net_8501), .D(net_3974), .SE(net_3884), .CK(net_10817) );
CLKBUF_X2 inst_12375 ( .A(net_12222), .Z(net_12223) );
CLKBUF_X2 inst_9591 ( .A(net_9438), .Z(net_9439) );
CLKBUF_X2 inst_16447 ( .A(net_16294), .Z(net_16295) );
NAND3_X2 inst_3909 ( .ZN(net_5629), .A1(net_5558), .A3(net_5492), .A2(net_5358) );
CLKBUF_X2 inst_18296 ( .A(net_17131), .Z(net_18144) );
SDFF_X2 inst_1869 ( .D(net_7271), .SI(net_6928), .Q(net_6928), .SE(net_6281), .CK(net_14103) );
SDFF_X2 inst_897 ( .SI(net_8709), .Q(net_8709), .SE(net_6195), .D(net_3965), .CK(net_13026) );
NAND3_X2 inst_3945 ( .A3(net_4468), .ZN(net_4467), .A1(net_4404), .A2(net_1679) );
CLKBUF_X2 inst_15592 ( .A(net_15439), .Z(net_15440) );
SDFF_X2 inst_1201 ( .D(net_7300), .SI(net_6877), .Q(net_6877), .SE(net_6282), .CK(net_15921) );
CLKBUF_X2 inst_11656 ( .A(net_11503), .Z(net_11504) );
AOI221_X2 inst_8760 ( .C2(net_6130), .B2(net_5535), .ZN(net_5472), .A(net_4952), .C1(net_1403), .B1(net_466) );
INV_X4 inst_5899 ( .A(net_6302), .ZN(net_2744) );
CLKBUF_X2 inst_9294 ( .A(net_9141), .Z(net_9142) );
CLKBUF_X2 inst_18331 ( .A(net_11425), .Z(net_18179) );
SDFF_X2 inst_1927 ( .SI(net_8054), .Q(net_8054), .D(net_2584), .SE(net_2508), .CK(net_18841) );
XNOR2_X2 inst_184 ( .ZN(net_1668), .B(net_1667), .A(net_1232) );
SDFF_X2 inst_1847 ( .D(net_7267), .SI(net_6884), .Q(net_6884), .SE(net_6284), .CK(net_16810) );
AOI21_X2 inst_8878 ( .B2(net_5871), .ZN(net_5867), .A(net_5861), .B1(net_2670) );
CLKBUF_X2 inst_12270 ( .A(net_11356), .Z(net_12118) );
CLKBUF_X2 inst_16312 ( .A(net_14953), .Z(net_16160) );
DFFS_X1 inst_6921 ( .D(net_6145), .CK(net_13661), .SN(x6501), .Q(x789) );
AOI221_X2 inst_8775 ( .B2(net_8236), .B1(net_5268), .C2(net_5267), .ZN(net_5264), .A(net_4914), .C1(net_173) );
AOI22_X2 inst_7742 ( .B1(net_6971), .A1(net_6931), .A2(net_5443), .B2(net_5442), .ZN(net_5438) );
CLKBUF_X2 inst_9409 ( .A(net_9256), .Z(net_9257) );
AND2_X4 inst_9125 ( .ZN(net_1403), .A2(net_920), .A1(net_177) );
CLKBUF_X2 inst_10919 ( .A(net_10766), .Z(net_10767) );
CLKBUF_X2 inst_15950 ( .A(net_15797), .Z(net_15798) );
CLKBUF_X2 inst_17270 ( .A(net_17117), .Z(net_17118) );
CLKBUF_X2 inst_17654 ( .A(net_17501), .Z(net_17502) );
SDFFR_X2 inst_2114 ( .QN(net_8908), .SE(net_6144), .D(net_5030), .SI(net_5029), .CK(net_17584), .RN(x6501) );
SDFFR_X1 inst_2784 ( .D(net_7379), .Q(net_7276), .SI(net_1941), .SE(net_1327), .CK(net_14770), .RN(x6501) );
INV_X2 inst_6330 ( .A(net_3179), .ZN(net_3119) );
CLKBUF_X2 inst_13817 ( .A(net_13664), .Z(net_13665) );
CLKBUF_X2 inst_13001 ( .A(net_12848), .Z(net_12849) );
CLKBUF_X2 inst_16105 ( .A(net_15952), .Z(net_15953) );
AND4_X2 inst_9036 ( .A3(net_4320), .ZN(net_2942), .A4(net_2769), .A2(net_2049), .A1(net_1872) );
CLKBUF_X2 inst_10538 ( .A(net_9281), .Z(net_10386) );
DFFR_X2 inst_7149 ( .QN(net_8950), .D(net_2891), .CK(net_14485), .RN(x6501) );
CLKBUF_X2 inst_16627 ( .A(net_16474), .Z(net_16475) );
CLKBUF_X2 inst_13458 ( .A(net_13305), .Z(net_13306) );
CLKBUF_X2 inst_13697 ( .A(net_10922), .Z(net_13545) );
NAND2_X2 inst_4377 ( .A1(net_7156), .A2(net_5166), .ZN(net_5080) );
NAND2_X2 inst_4301 ( .A1(net_7052), .A2(net_5162), .ZN(net_5156) );
CLKBUF_X2 inst_16046 ( .A(net_13667), .Z(net_15894) );
CLKBUF_X2 inst_13432 ( .A(net_13279), .Z(net_13280) );
AOI22_X2 inst_8537 ( .B1(net_6725), .A1(net_6692), .B2(net_6202), .A2(net_3520), .ZN(net_3403) );
CLKBUF_X2 inst_16188 ( .A(net_15590), .Z(net_16036) );
CLKBUF_X2 inst_15018 ( .A(net_14865), .Z(net_14866) );
INV_X4 inst_5106 ( .ZN(net_5688), .A(net_5597) );
SDFF_X2 inst_1410 ( .SI(net_7267), .Q(net_7084), .D(net_7084), .SE(net_6278), .CK(net_16866) );
CLKBUF_X2 inst_14943 ( .A(net_14790), .Z(net_14791) );
CLKBUF_X2 inst_10675 ( .A(net_10522), .Z(net_10523) );
CLKBUF_X2 inst_16510 ( .A(net_16357), .Z(net_16358) );
NAND2_X2 inst_4424 ( .A1(net_6862), .A2(net_5016), .ZN(net_5003) );
DFFR_X2 inst_7028 ( .QN(net_9011), .D(net_5689), .CK(net_11167), .RN(x6501) );
INV_X4 inst_5994 ( .ZN(net_918), .A(net_400) );
CLKBUF_X2 inst_19067 ( .A(net_17612), .Z(net_18915) );
CLKBUF_X2 inst_10210 ( .A(net_10057), .Z(net_10058) );
CLKBUF_X2 inst_18952 ( .A(net_18799), .Z(net_18800) );
INV_X1 inst_6653 ( .A(net_7414), .ZN(net_569) );
CLKBUF_X2 inst_18284 ( .A(net_18131), .Z(net_18132) );
SDFFS_X2 inst_2074 ( .SI(net_7387), .SE(net_2795), .Q(net_176), .D(net_176), .CK(net_14666), .SN(x6501) );
CLKBUF_X2 inst_11330 ( .A(net_11177), .Z(net_11178) );
DFFR_X2 inst_7296 ( .QN(net_8947), .D(net_1371), .CK(net_16285), .RN(x6501) );
NAND2_X2 inst_4823 ( .ZN(net_1166), .A2(net_863), .A1(net_180) );
SDFF_X2 inst_1236 ( .Q(net_7814), .D(net_7814), .SE(net_2730), .SI(net_2702), .CK(net_18093) );
XNOR2_X2 inst_221 ( .B(net_6821), .ZN(net_1394), .A(net_1393) );
INV_X4 inst_5112 ( .A(net_5272), .ZN(net_4938) );
INV_X4 inst_5929 ( .A(net_6368), .ZN(net_1241) );
NOR3_X2 inst_3313 ( .A3(net_7502), .A2(net_7501), .ZN(net_1436), .A1(net_1435) );
CLKBUF_X2 inst_12640 ( .A(net_12487), .Z(net_12488) );
NOR2_X2 inst_3562 ( .ZN(net_1727), .A2(net_1622), .A1(net_602) );
CLKBUF_X2 inst_9545 ( .A(net_9392), .Z(net_9393) );
CLKBUF_X2 inst_13502 ( .A(net_13349), .Z(net_13350) );
CLKBUF_X2 inst_18635 ( .A(net_18482), .Z(net_18483) );
SDFFR_X2 inst_2334 ( .QN(net_6347), .SI(net_2760), .D(net_2739), .SE(net_2320), .CK(net_17819), .RN(x6501) );
CLKBUF_X2 inst_11967 ( .A(net_11814), .Z(net_11815) );
CLKBUF_X2 inst_17261 ( .A(net_17108), .Z(net_17109) );
SDFFR_X2 inst_2210 ( .Q(net_7444), .D(net_7444), .SE(net_2863), .CK(net_12821), .SI(x13626), .RN(x6501) );
INV_X4 inst_6040 ( .A(net_7489), .ZN(net_4890) );
INV_X8 inst_5028 ( .ZN(net_3884), .A(net_3303) );
SDFFR_X2 inst_2590 ( .D(net_7388), .QN(net_7248), .SI(net_1946), .SE(net_1379), .CK(net_18108), .RN(x6501) );
CLKBUF_X2 inst_11577 ( .A(net_11424), .Z(net_11425) );
CLKBUF_X2 inst_10949 ( .A(net_10285), .Z(net_10797) );
CLKBUF_X2 inst_10435 ( .A(net_9714), .Z(net_10283) );
INV_X8 inst_5025 ( .ZN(net_3983), .A(net_3321) );
CLKBUF_X2 inst_16947 ( .A(net_16794), .Z(net_16795) );
CLKBUF_X2 inst_18739 ( .A(net_18586), .Z(net_18587) );
CLKBUF_X2 inst_13341 ( .A(net_9677), .Z(net_13189) );
CLKBUF_X2 inst_18340 ( .A(net_18187), .Z(net_18188) );
CLKBUF_X2 inst_17900 ( .A(net_17747), .Z(net_17748) );
CLKBUF_X2 inst_12451 ( .A(net_10325), .Z(net_12299) );
NAND2_X2 inst_4459 ( .ZN(net_4933), .A2(net_4712), .A1(net_4494) );
CLKBUF_X2 inst_15261 ( .A(net_15108), .Z(net_15109) );
CLKBUF_X2 inst_14028 ( .A(net_13875), .Z(net_13876) );
SDFF_X2 inst_1117 ( .D(net_7321), .SI(net_6563), .Q(net_6563), .SE(net_3070), .CK(net_9150) );
DFFR_X2 inst_7343 ( .Q(net_7337), .CK(net_11712), .D(x12940), .RN(x6501) );
NAND2_X4 inst_4015 ( .ZN(net_4455), .A1(net_4374), .A2(net_4359) );
CLKBUF_X2 inst_11374 ( .A(net_11221), .Z(net_11222) );
CLKBUF_X2 inst_13909 ( .A(net_13756), .Z(net_13757) );
DFFS_X2 inst_6887 ( .QN(net_6113), .D(net_2944), .CK(net_14471), .SN(x6501) );
SDFFR_X1 inst_2725 ( .SI(net_9037), .Q(net_9037), .D(net_7466), .SE(net_3208), .CK(net_10662), .RN(x6501) );
HA_X1 inst_6681 ( .S(net_3043), .CO(net_3042), .B(net_2875), .A(x2693) );
INV_X4 inst_5141 ( .ZN(net_3889), .A(net_3598) );
CLKBUF_X2 inst_14476 ( .A(net_11208), .Z(net_14324) );
AOI22_X2 inst_8204 ( .A1(net_8608), .B1(net_8423), .A2(net_3864), .B2(net_3863), .ZN(net_3832) );
SDFF_X2 inst_1610 ( .Q(net_8116), .D(net_8116), .SI(net_2709), .SE(net_2541), .CK(net_15766) );
XNOR2_X2 inst_334 ( .B(net_7392), .A(net_6374), .ZN(net_793) );
CLKBUF_X2 inst_13337 ( .A(net_13184), .Z(net_13185) );
SDFF_X2 inst_1042 ( .SI(net_7333), .Q(net_6707), .D(net_6707), .SE(net_3125), .CK(net_9426) );
CLKBUF_X2 inst_14190 ( .A(net_14037), .Z(net_14038) );
INV_X4 inst_5961 ( .A(net_7478), .ZN(net_3128) );
CLKBUF_X2 inst_15850 ( .A(net_14182), .Z(net_15698) );
INV_X4 inst_5595 ( .A(net_6458), .ZN(net_3032) );
AOI22_X2 inst_8153 ( .B1(net_8121), .A1(net_7883), .A2(net_6098), .ZN(net_6054), .B2(net_4190) );
CLKBUF_X2 inst_17068 ( .A(net_15005), .Z(net_16916) );
CLKBUF_X2 inst_18497 ( .A(net_18344), .Z(net_18345) );
AOI22_X2 inst_8058 ( .B1(net_8207), .A1(net_7697), .B2(net_6099), .A2(net_4399), .ZN(net_4084) );
SDFF_X2 inst_595 ( .SI(net_8387), .Q(net_8387), .SE(net_3969), .D(net_3944), .CK(net_10840) );
CLKBUF_X2 inst_13255 ( .A(net_13102), .Z(net_13103) );
MUX2_X2 inst_5002 ( .A(net_9019), .Z(net_3938), .B(net_1444), .S(net_622) );
AOI22_X2 inst_8222 ( .B1(net_8869), .A1(net_8314), .B2(net_6252), .A2(net_4345), .ZN(net_3814) );
INV_X2 inst_6343 ( .ZN(net_2527), .A(net_2486) );
CLKBUF_X2 inst_13554 ( .A(net_13401), .Z(net_13402) );
AOI211_X2 inst_9014 ( .C2(net_5463), .A(net_4834), .ZN(net_4833), .B(net_4560), .C1(net_2555) );
CLKBUF_X2 inst_19035 ( .A(net_15437), .Z(net_18883) );
NAND2_X2 inst_4688 ( .ZN(net_6216), .A2(net_6157), .A1(net_1460) );
CLKBUF_X2 inst_12658 ( .A(net_12505), .Z(net_12506) );
CLKBUF_X2 inst_15451 ( .A(net_15298), .Z(net_15299) );
CLKBUF_X2 inst_17833 ( .A(net_17680), .Z(net_17681) );
CLKBUF_X2 inst_17219 ( .A(net_17066), .Z(net_17067) );
NAND2_X2 inst_4798 ( .ZN(net_3278), .A2(net_1378), .A1(net_1150) );
NAND4_X2 inst_3849 ( .A4(net_7210), .ZN(net_1624), .A2(net_1617), .A3(net_1477), .A1(net_1279) );
CLKBUF_X2 inst_12205 ( .A(net_9444), .Z(net_12053) );
CLKBUF_X2 inst_15575 ( .A(net_15422), .Z(net_15423) );
CLKBUF_X2 inst_15840 ( .A(net_15687), .Z(net_15688) );
CLKBUF_X2 inst_19188 ( .A(net_11432), .Z(net_19036) );
SDFF_X2 inst_1029 ( .SI(net_7334), .Q(net_6741), .D(net_6741), .SE(net_3124), .CK(net_12017) );
INV_X4 inst_5413 ( .ZN(net_1087), .A(net_867) );
HA_X1 inst_6666 ( .S(net_3268), .CO(net_3267), .B(net_3103), .A(x2908) );
CLKBUF_X2 inst_9246 ( .A(net_9093), .Z(net_9094) );
DFF_X1 inst_6841 ( .Q(net_6431), .D(net_3606), .CK(net_17972) );
DFFR_X2 inst_7032 ( .QN(net_7490), .D(net_5042), .CK(net_16593), .RN(x6501) );
INV_X2 inst_6245 ( .ZN(net_4861), .A(net_4756) );
INV_X2 inst_6551 ( .A(net_6376), .ZN(net_2120) );
INV_X4 inst_5767 ( .A(net_6367), .ZN(net_558) );
CLKBUF_X2 inst_13048 ( .A(net_12319), .Z(net_12896) );
CLKBUF_X2 inst_10067 ( .A(net_9914), .Z(net_9915) );
INV_X2 inst_6443 ( .A(net_1241), .ZN(net_614) );
CLKBUF_X2 inst_14404 ( .A(net_14251), .Z(net_14252) );
SDFF_X2 inst_1534 ( .Q(net_7883), .D(net_7883), .SI(net_2573), .SE(net_2543), .CK(net_15277) );
CLKBUF_X2 inst_9985 ( .A(net_9594), .Z(net_9833) );
XNOR2_X2 inst_319 ( .A(net_1780), .ZN(net_944), .B(net_943) );
AND2_X4 inst_9108 ( .ZN(net_2122), .A1(net_1936), .A2(net_1935) );
SDFFR_X2 inst_2422 ( .QN(net_9007), .D(net_2680), .SI(net_2427), .SE(net_2266), .CK(net_16251), .RN(x6501) );
CLKBUF_X2 inst_12745 ( .A(net_12592), .Z(net_12593) );
CLKBUF_X2 inst_10688 ( .A(net_10407), .Z(net_10536) );
SDFF_X2 inst_649 ( .Q(net_8420), .D(net_8420), .SI(net_3945), .SE(net_3934), .CK(net_13045) );
CLKBUF_X2 inst_18724 ( .A(net_9835), .Z(net_18572) );
INV_X4 inst_5790 ( .A(net_7215), .ZN(net_692) );
CLKBUF_X2 inst_18676 ( .A(net_18523), .Z(net_18524) );
CLKBUF_X2 inst_15166 ( .A(net_15013), .Z(net_15014) );
SDFFR_X2 inst_2597 ( .D(net_7396), .QN(net_7256), .SI(net_1939), .SE(net_1379), .CK(net_18314), .RN(x6501) );
AOI22_X2 inst_8504 ( .B1(net_6549), .A1(net_6516), .A2(net_6137), .B2(net_6104), .ZN(net_3436) );
CLKBUF_X2 inst_16379 ( .A(net_16226), .Z(net_16227) );
CLKBUF_X2 inst_14269 ( .A(net_14116), .Z(net_14117) );
INV_X4 inst_5569 ( .A(net_7343), .ZN(net_2185) );
INV_X4 inst_5185 ( .ZN(net_2881), .A(net_2834) );
CLKBUF_X2 inst_12227 ( .A(net_12074), .Z(net_12075) );
INV_X4 inst_6059 ( .ZN(net_494), .A(x352) );
SDFF_X2 inst_1575 ( .Q(net_8025), .D(net_8025), .SI(net_2576), .SE(net_2545), .CK(net_16047) );
CLKBUF_X2 inst_17453 ( .A(net_17300), .Z(net_17301) );
CLKBUF_X2 inst_9644 ( .A(net_9491), .Z(net_9492) );
CLKBUF_X2 inst_16300 ( .A(net_16147), .Z(net_16148) );
INV_X4 inst_5522 ( .ZN(net_670), .A(net_669) );
SDFF_X2 inst_1258 ( .Q(net_8097), .D(net_8097), .SI(net_2722), .SE(net_2707), .CK(net_18815) );
OAI21_X2 inst_3141 ( .B2(net_2060), .ZN(net_2055), .A(net_2054), .B1(net_1523) );
CLKBUF_X2 inst_10148 ( .A(net_9995), .Z(net_9996) );
NAND3_X2 inst_3921 ( .ZN(net_5617), .A1(net_5546), .A3(net_5480), .A2(net_5307) );
CLKBUF_X2 inst_16820 ( .A(net_16667), .Z(net_16668) );
SDFF_X2 inst_1957 ( .D(net_7298), .SI(net_7035), .Q(net_7035), .SE(net_6277), .CK(net_18176) );
INV_X4 inst_5151 ( .ZN(net_3231), .A(net_3188) );
CLKBUF_X2 inst_9524 ( .A(net_9371), .Z(net_9372) );
CLKBUF_X2 inst_13860 ( .A(net_13707), .Z(net_13708) );
DFFR_X1 inst_7446 ( .QN(net_8926), .D(net_4757), .CK(net_13967), .RN(x6501) );
CLKBUF_X2 inst_10456 ( .A(net_10154), .Z(net_10304) );
CLKBUF_X2 inst_13813 ( .A(net_12825), .Z(net_13661) );
NAND2_X2 inst_4624 ( .A2(net_6144), .ZN(net_2593), .A1(net_2592) );
AOI22_X2 inst_7811 ( .A2(net_8238), .B2(net_6144), .A1(net_4764), .ZN(net_4753), .B1(net_4518) );
CLKBUF_X2 inst_12458 ( .A(net_12305), .Z(net_12306) );
CLKBUF_X2 inst_11257 ( .A(net_11104), .Z(net_11105) );
CLKBUF_X2 inst_18597 ( .A(net_18444), .Z(net_18445) );
INV_X4 inst_6062 ( .A(net_6471), .ZN(net_1542) );
CLKBUF_X2 inst_9254 ( .A(net_9101), .Z(net_9102) );
DFFR_X1 inst_7428 ( .QN(net_8929), .D(net_4859), .CK(net_16697), .RN(x6501) );
AOI22_X2 inst_7778 ( .B1(net_6968), .A1(net_6928), .A2(net_5443), .B2(net_5442), .ZN(net_5291) );
INV_X2 inst_6608 ( .A(net_6185), .ZN(net_6184) );
OAI21_X2 inst_2983 ( .B1(net_7630), .ZN(net_5929), .A(net_5853), .B2(net_5852) );
DFFR_X1 inst_7421 ( .QN(net_7514), .D(net_4939), .CK(net_14862), .RN(x6501) );
CLKBUF_X2 inst_13233 ( .A(net_13080), .Z(net_13081) );
CLKBUF_X2 inst_13584 ( .A(net_10130), .Z(net_13432) );
AOI221_X2 inst_8862 ( .C1(net_8901), .B2(net_6160), .ZN(net_4729), .A(net_1887), .C2(net_1886), .B1(net_878) );
CLKBUF_X2 inst_9969 ( .A(net_9672), .Z(net_9817) );
CLKBUF_X2 inst_12881 ( .A(net_12728), .Z(net_12729) );
SDFF_X2 inst_1120 ( .D(net_7325), .SI(net_6567), .Q(net_6567), .SE(net_3070), .CK(net_9125) );
INV_X2 inst_6238 ( .ZN(net_5281), .A(net_5032) );
CLKBUF_X2 inst_12986 ( .A(net_12833), .Z(net_12834) );
CLKBUF_X2 inst_16035 ( .A(net_15882), .Z(net_15883) );
AOI22_X2 inst_8545 ( .B1(net_6727), .A1(net_6694), .B2(net_6202), .A2(net_3520), .ZN(net_3395) );
CLKBUF_X2 inst_15029 ( .A(net_14876), .Z(net_14877) );
OAI211_X2 inst_3184 ( .ZN(net_5525), .C2(net_5036), .B(net_4731), .A(net_1590), .C1(net_1068) );
INV_X2 inst_6398 ( .ZN(net_1161), .A(net_1160) );
CLKBUF_X2 inst_9715 ( .A(net_9562), .Z(net_9563) );
SDFF_X2 inst_947 ( .SI(net_7330), .Q(net_6704), .D(net_6704), .SE(net_3125), .CK(net_11336) );
SDFF_X2 inst_731 ( .SI(net_8340), .Q(net_8340), .D(net_3947), .SE(net_3880), .CK(net_12433) );
CLKBUF_X2 inst_15381 ( .A(net_13937), .Z(net_15229) );
CLKBUF_X2 inst_10909 ( .A(net_9501), .Z(net_10757) );
CLKBUF_X2 inst_13788 ( .A(net_13635), .Z(net_13636) );
CLKBUF_X2 inst_15005 ( .A(net_14852), .Z(net_14853) );
SDFFR_X2 inst_2459 ( .SI(net_7375), .SE(net_2723), .D(net_2641), .QN(net_156), .CK(net_17807), .RN(x6501) );
DFFR_X2 inst_7165 ( .QN(net_8945), .D(net_2651), .CK(net_16310), .RN(x6501) );
XNOR2_X2 inst_301 ( .ZN(net_979), .A(net_978), .B(net_191) );
SDFF_X2 inst_363 ( .SI(net_8327), .Q(net_8327), .SE(net_3978), .D(net_3940), .CK(net_10306) );
SDFFR_X2 inst_2141 ( .SI(net_7204), .Q(net_7204), .D(net_6455), .SE(net_4362), .CK(net_14560), .RN(x6501) );
CLKBUF_X2 inst_12041 ( .A(net_11036), .Z(net_11889) );
INV_X2 inst_6609 ( .A(net_6186), .ZN(net_6185) );
DFFR_X2 inst_7079 ( .QN(net_7648), .D(net_3897), .CK(net_12691), .RN(x6501) );
CLKBUF_X2 inst_13213 ( .A(net_12254), .Z(net_13061) );
AOI22_X2 inst_7870 ( .B2(net_5609), .A2(net_5267), .ZN(net_4571), .B1(net_361), .A1(net_165) );
CLKBUF_X2 inst_14021 ( .A(net_13868), .Z(net_13869) );
CLKBUF_X2 inst_19000 ( .A(net_10037), .Z(net_18848) );
NAND2_X2 inst_4706 ( .ZN(net_1860), .A2(net_1771), .A1(net_1330) );
NAND2_X2 inst_4348 ( .A1(net_7107), .A2(net_5164), .ZN(net_5109) );
NAND4_X2 inst_3729 ( .ZN(net_4301), .A1(net_4142), .A2(net_4141), .A3(net_4140), .A4(net_4139) );
CLKBUF_X2 inst_14312 ( .A(net_10525), .Z(net_14160) );
AOI22_X2 inst_8521 ( .B1(net_6721), .A1(net_6688), .B2(net_6202), .A2(net_3520), .ZN(net_3419) );
DFFR_X1 inst_7548 ( .Q(net_7628), .D(net_915), .CK(net_15710), .RN(x6501) );
CLKBUF_X2 inst_10430 ( .A(net_9394), .Z(net_10278) );
AOI22_X2 inst_8345 ( .B1(net_8700), .A1(net_8663), .B2(net_6109), .A2(net_3857), .ZN(net_3702) );
CLKBUF_X2 inst_9282 ( .A(net_9129), .Z(net_9130) );
SDFFR_X1 inst_2650 ( .D(net_6773), .SE(net_4506), .CK(net_9198), .RN(x6501), .SI(x1690), .Q(x1690) );
CLKBUF_X2 inst_11687 ( .A(net_11534), .Z(net_11535) );
CLKBUF_X2 inst_14559 ( .A(net_12473), .Z(net_14407) );
CLKBUF_X2 inst_16102 ( .A(net_10856), .Z(net_15950) );
NAND2_X2 inst_4508 ( .A1(net_8965), .A2(net_6206), .ZN(net_4387) );
CLKBUF_X2 inst_16791 ( .A(net_16638), .Z(net_16639) );
AOI22_X2 inst_7943 ( .B1(net_8021), .A1(net_7987), .B2(net_6102), .A2(net_6097), .ZN(net_4182) );
CLKBUF_X2 inst_16134 ( .A(net_15981), .Z(net_15982) );
CLKBUF_X2 inst_11626 ( .A(net_11473), .Z(net_11474) );
CLKBUF_X2 inst_9490 ( .A(net_9337), .Z(net_9338) );
CLKBUF_X2 inst_11666 ( .A(net_11513), .Z(net_11514) );
CLKBUF_X2 inst_18315 ( .A(net_18162), .Z(net_18163) );
OAI211_X2 inst_3189 ( .ZN(net_4819), .A(net_4672), .B(net_4476), .C2(net_4370), .C1(net_1903) );
AOI21_X2 inst_8918 ( .ZN(net_5752), .A(net_5745), .B2(net_5593), .B1(net_4788) );
CLKBUF_X2 inst_12818 ( .A(net_12665), .Z(net_12666) );
DFF_X1 inst_6855 ( .Q(net_6443), .D(net_3626), .CK(net_17890) );
INV_X4 inst_5985 ( .A(net_8970), .ZN(net_677) );
INV_X4 inst_5548 ( .ZN(net_1060), .A(net_638) );
CLKBUF_X2 inst_14188 ( .A(net_14035), .Z(net_14036) );
CLKBUF_X2 inst_10902 ( .A(net_9101), .Z(net_10750) );
SDFF_X2 inst_684 ( .Q(net_8681), .D(net_8681), .SI(net_3959), .SE(net_3935), .CK(net_13189) );
INV_X2 inst_6263 ( .A(net_8242), .ZN(net_4634) );
NAND2_X2 inst_4400 ( .A1(net_7046), .A2(net_5162), .ZN(net_5057) );
OAI211_X2 inst_3177 ( .B(net_6792), .A(net_6185), .C2(net_6146), .ZN(net_5838), .C1(net_1898) );
CLKBUF_X2 inst_12187 ( .A(net_12034), .Z(net_12035) );
MUX2_X2 inst_4930 ( .A(net_8261), .Z(net_3120), .S(net_2996), .B(net_1697) );
CLKBUF_X2 inst_10437 ( .A(net_10284), .Z(net_10285) );
AOI22_X2 inst_7965 ( .A1(net_7956), .B1(net_7786), .A2(net_6092), .B2(net_6091), .ZN(net_4163) );
CLKBUF_X2 inst_18585 ( .A(net_18432), .Z(net_18433) );
CLKBUF_X2 inst_11857 ( .A(net_11704), .Z(net_11705) );
SDFF_X2 inst_1138 ( .D(net_7317), .SI(net_6559), .Q(net_6559), .SE(net_3070), .CK(net_11996) );
INV_X2 inst_6568 ( .A(net_6360), .ZN(net_2131) );
SDFF_X2 inst_1004 ( .D(net_7315), .SI(net_6623), .Q(net_6623), .SE(net_3123), .CK(net_9939) );
XNOR2_X2 inst_189 ( .ZN(net_1603), .B(net_1119), .A(net_932) );
CLKBUF_X2 inst_9316 ( .A(net_9163), .Z(net_9164) );
SDFFR_X2 inst_2450 ( .D(net_3272), .SE(net_2313), .SI(net_418), .Q(net_418), .CK(net_16655), .RN(x6501) );
CLKBUF_X2 inst_13248 ( .A(net_13095), .Z(net_13096) );
DFFR_X1 inst_7437 ( .QN(net_8917), .D(net_4846), .CK(net_16688), .RN(x6501) );
AOI222_X1 inst_8597 ( .B2(net_6775), .B1(net_5835), .C2(net_5832), .A2(net_5830), .ZN(net_5829), .A1(net_2979), .C1(x2805) );
CLKBUF_X2 inst_16190 ( .A(net_13850), .Z(net_16038) );
DFFR_X1 inst_7430 ( .QN(net_8937), .D(net_4857), .CK(net_14596), .RN(x6501) );
XOR2_X2 inst_62 ( .Z(net_932), .A(net_931), .B(net_930) );
CLKBUF_X2 inst_9529 ( .A(net_9376), .Z(net_9377) );
CLKBUF_X2 inst_11006 ( .A(net_10853), .Z(net_10854) );
NAND2_X2 inst_4696 ( .A2(net_6162), .ZN(net_2090), .A1(net_829) );
NAND4_X2 inst_3743 ( .ZN(net_4287), .A1(net_4058), .A2(net_4057), .A3(net_4056), .A4(net_4055) );
CLKBUF_X2 inst_16247 ( .A(net_16094), .Z(net_16095) );
OR2_X4 inst_2860 ( .ZN(net_6281), .A2(net_2199), .A1(net_1922) );
INV_X4 inst_5194 ( .ZN(net_4922), .A(net_2642) );
CLKBUF_X2 inst_17713 ( .A(net_17560), .Z(net_17561) );
AOI22_X2 inst_8387 ( .B1(net_8672), .A1(net_8635), .B2(net_6109), .A2(net_3857), .ZN(net_3661) );
CLKBUF_X2 inst_14496 ( .A(net_11793), .Z(net_14344) );
INV_X4 inst_5888 ( .A(net_5956), .ZN(net_1106) );
CLKBUF_X2 inst_11266 ( .A(net_9238), .Z(net_11114) );
CLKBUF_X2 inst_17344 ( .A(net_17191), .Z(net_17192) );
CLKBUF_X2 inst_11162 ( .A(net_9623), .Z(net_11010) );
CLKBUF_X2 inst_13956 ( .A(net_13803), .Z(net_13804) );
DFFR_X2 inst_7344 ( .Q(net_7311), .CK(net_11383), .D(x13185), .RN(x6501) );
AOI22_X2 inst_8252 ( .B1(net_8725), .A1(net_8503), .ZN(net_6065), .B2(net_4350), .A2(net_4349) );
CLKBUF_X2 inst_12416 ( .A(net_12263), .Z(net_12264) );
NAND2_X2 inst_4482 ( .A2(net_5267), .ZN(net_4496), .A1(net_167) );
CLKBUF_X2 inst_15462 ( .A(net_15309), .Z(net_15310) );
CLKBUF_X2 inst_16713 ( .A(net_16560), .Z(net_16561) );
AOI22_X2 inst_7903 ( .B1(net_7191), .A2(net_6442), .B2(net_5655), .A1(net_5654), .ZN(net_4524) );
CLKBUF_X2 inst_18051 ( .A(net_11977), .Z(net_17899) );
SDFF_X2 inst_791 ( .SI(net_8362), .Q(net_8362), .D(net_3953), .SE(net_3880), .CK(net_10238) );
CLKBUF_X2 inst_18016 ( .A(net_17863), .Z(net_17864) );
CLKBUF_X2 inst_10427 ( .A(net_10274), .Z(net_10275) );
CLKBUF_X2 inst_13371 ( .A(net_13218), .Z(net_13219) );
SDFF_X2 inst_2021 ( .SI(net_7928), .Q(net_7928), .D(net_2718), .SE(net_2461), .CK(net_18345) );
CLKBUF_X2 inst_9631 ( .A(net_9478), .Z(net_9479) );
CLKBUF_X2 inst_18424 ( .A(net_18271), .Z(net_18272) );
NAND2_X2 inst_4379 ( .A1(net_7076), .A2(net_5162), .ZN(net_5078) );
INV_X4 inst_5668 ( .A(net_7477), .ZN(net_3129) );
CLKBUF_X2 inst_13326 ( .A(net_13173), .Z(net_13174) );
INV_X4 inst_5086 ( .ZN(net_5728), .A(net_5701) );
CLKBUF_X2 inst_15107 ( .A(net_12766), .Z(net_14955) );
CLKBUF_X2 inst_12811 ( .A(net_12658), .Z(net_12659) );
CLKBUF_X2 inst_17983 ( .A(net_17830), .Z(net_17831) );
CLKBUF_X2 inst_14670 ( .A(net_14517), .Z(net_14518) );
AOI22_X2 inst_8576 ( .B2(net_7169), .A2(net_7168), .A1(net_1830), .B1(net_1829), .ZN(net_1652) );
CLKBUF_X2 inst_14399 ( .A(net_13426), .Z(net_14247) );
CLKBUF_X2 inst_11924 ( .A(net_11771), .Z(net_11772) );
CLKBUF_X2 inst_13020 ( .A(net_12867), .Z(net_12868) );
CLKBUF_X2 inst_11888 ( .A(net_11735), .Z(net_11736) );
AOI22_X2 inst_7848 ( .B2(net_5595), .A2(net_4809), .ZN(net_4660), .A1(net_723), .B1(net_317) );
AOI22_X2 inst_8142 ( .A1(net_7949), .B1(net_7779), .A2(net_6092), .B2(net_6091), .ZN(net_4009) );
INV_X4 inst_6143 ( .A(net_6133), .ZN(net_6129) );
DFFR_X2 inst_7304 ( .D(net_7641), .QN(net_7638), .CK(net_15653), .RN(x6501) );
CLKBUF_X2 inst_12864 ( .A(net_12614), .Z(net_12712) );
NAND2_X2 inst_4404 ( .A1(net_7128), .A2(net_5166), .ZN(net_5053) );
AOI21_X2 inst_8937 ( .B2(net_5871), .ZN(net_5665), .A(net_5664), .B1(net_2686) );
CLKBUF_X2 inst_18119 ( .A(net_17966), .Z(net_17967) );
AND2_X4 inst_9054 ( .A2(net_3356), .ZN(net_3353), .A1(net_3320) );
AOI22_X2 inst_8154 ( .B1(net_8189), .A1(net_7679), .B2(net_6099), .A2(net_4399), .ZN(net_3998) );
INV_X2 inst_6581 ( .A(net_7669), .ZN(net_919) );
CLKBUF_X2 inst_17651 ( .A(net_14767), .Z(net_17499) );
CLKBUF_X2 inst_11261 ( .A(net_11108), .Z(net_11109) );
CLKBUF_X2 inst_16130 ( .A(net_15977), .Z(net_15978) );
CLKBUF_X2 inst_18395 ( .A(net_18242), .Z(net_18243) );
DFF_X1 inst_6716 ( .QN(net_6793), .D(net_5620), .CK(net_11596) );
CLKBUF_X2 inst_15046 ( .A(net_14893), .Z(net_14894) );
INV_X4 inst_5541 ( .A(net_1855), .ZN(net_649) );
NAND2_X4 inst_4018 ( .A1(net_6273), .ZN(net_4374), .A2(net_4373) );
CLKBUF_X2 inst_16430 ( .A(net_16277), .Z(net_16278) );
INV_X4 inst_5636 ( .A(net_6315), .ZN(net_2725) );
SDFFR_X2 inst_2219 ( .Q(net_7453), .D(net_7453), .SE(net_2863), .CK(net_12923), .SI(x13553), .RN(x6501) );
CLKBUF_X2 inst_17854 ( .A(net_11666), .Z(net_17702) );
AOI22_X2 inst_8331 ( .B1(net_8698), .A1(net_8661), .B2(net_6109), .A2(net_3857), .ZN(net_3715) );
AOI21_X2 inst_8884 ( .B2(net_5871), .ZN(net_5839), .A(net_5795), .B1(x225) );
SDFF_X2 inst_1284 ( .Q(net_7833), .D(net_7833), .SE(net_2730), .SI(net_2639), .CK(net_17156) );
SDFF_X2 inst_546 ( .Q(net_8690), .D(net_8690), .SI(net_3942), .SE(net_3935), .CK(net_10566) );
CLKBUF_X2 inst_18970 ( .A(net_18817), .Z(net_18818) );
SDFFR_X2 inst_2465 ( .SE(net_2260), .Q(net_308), .D(net_308), .CK(net_10398), .RN(x6501), .SI(x3604) );
SDFF_X2 inst_704 ( .SI(net_8602), .Q(net_8602), .SE(net_3984), .D(net_3946), .CK(net_10750) );
CLKBUF_X2 inst_9301 ( .A(net_9148), .Z(net_9149) );
CLKBUF_X2 inst_16128 ( .A(net_15975), .Z(net_15976) );
NAND2_X2 inst_4542 ( .ZN(net_3357), .A2(net_3356), .A1(net_3326) );
DFFR_X2 inst_7084 ( .QN(net_7650), .D(net_3891), .CK(net_12676), .RN(x6501) );
INV_X4 inst_5558 ( .ZN(net_629), .A(net_628) );
AOI22_X2 inst_8285 ( .B1(net_8582), .A1(net_8471), .A2(net_6263), .B2(net_6262), .ZN(net_3757) );
SDFFR_X2 inst_2226 ( .Q(net_7446), .D(net_7446), .SE(net_2863), .CK(net_12808), .SI(x13612), .RN(x6501) );
CLKBUF_X2 inst_15538 ( .A(net_15385), .Z(net_15386) );
INV_X4 inst_5467 ( .ZN(net_817), .A(net_754) );
CLKBUF_X2 inst_17113 ( .A(net_16960), .Z(net_16961) );
CLKBUF_X2 inst_18915 ( .A(net_13625), .Z(net_18763) );
CLKBUF_X2 inst_17299 ( .A(net_17146), .Z(net_17147) );
CLKBUF_X2 inst_16652 ( .A(net_16499), .Z(net_16500) );
CLKBUF_X2 inst_17926 ( .A(net_17773), .Z(net_17774) );
DFFR_X2 inst_6986 ( .QN(net_6311), .D(net_5916), .CK(net_13960), .RN(x6501) );
CLKBUF_X2 inst_11476 ( .A(net_11323), .Z(net_11324) );
AOI21_X2 inst_8983 ( .ZN(net_1898), .A(net_1897), .B2(net_1629), .B1(net_962) );
CLKBUF_X2 inst_11523 ( .A(net_11370), .Z(net_11371) );
CLKBUF_X2 inst_17054 ( .A(net_16901), .Z(net_16902) );
CLKBUF_X2 inst_13885 ( .A(net_12481), .Z(net_13733) );
INV_X4 inst_5211 ( .ZN(net_2380), .A(net_2298) );
CLKBUF_X2 inst_11467 ( .A(net_11314), .Z(net_11315) );
SDFF_X2 inst_1342 ( .SI(net_7710), .Q(net_7710), .D(net_2708), .SE(net_2559), .CK(net_15537) );
OAI221_X2 inst_2971 ( .B2(net_2489), .ZN(net_2451), .C2(net_2450), .A(net_2271), .B1(net_1753), .C1(net_675) );
NAND2_X2 inst_4549 ( .A2(net_3367), .A1(net_3315), .ZN(net_3314) );
DFFR_X1 inst_7483 ( .QN(net_7428), .D(net_4206), .CK(net_12384), .RN(x6501) );
INV_X4 inst_6012 ( .A(net_7431), .ZN(net_3269) );
CLKBUF_X2 inst_10551 ( .A(net_9064), .Z(net_10399) );
NAND3_X2 inst_3933 ( .ZN(net_5517), .A1(net_5279), .A2(net_4657), .A3(net_4568) );
SDFF_X2 inst_1656 ( .SI(net_7711), .Q(net_7711), .D(net_2658), .SE(net_2559), .CK(net_15262) );
INV_X4 inst_5881 ( .A(net_8902), .ZN(net_1886) );
SDFF_X2 inst_1881 ( .D(net_7291), .SI(net_6988), .Q(net_6988), .SE(net_6283), .CK(net_15317) );
CLKBUF_X2 inst_18894 ( .A(net_18741), .Z(net_18742) );
CLKBUF_X2 inst_18729 ( .A(net_18576), .Z(net_18577) );
INV_X4 inst_5590 ( .A(net_7351), .ZN(net_2207) );
OAI21_X2 inst_3034 ( .B1(net_4850), .ZN(net_4848), .B2(net_4847), .A(net_2631) );
XNOR2_X2 inst_295 ( .A(net_1462), .ZN(net_987), .B(net_189) );
CLKBUF_X2 inst_15507 ( .A(net_15354), .Z(net_15355) );
CLKBUF_X2 inst_18812 ( .A(net_18659), .Z(net_18660) );
CLKBUF_X2 inst_17700 ( .A(net_9089), .Z(net_17548) );
CLKBUF_X2 inst_17665 ( .A(net_17512), .Z(net_17513) );
AOI21_X2 inst_8971 ( .ZN(net_6090), .B2(net_5986), .B1(net_2321), .A(net_1289) );
CLKBUF_X2 inst_13018 ( .A(net_12865), .Z(net_12866) );
SDFF_X2 inst_607 ( .SI(net_8401), .Q(net_8401), .SE(net_3969), .D(net_3940), .CK(net_10260) );
INV_X2 inst_6484 ( .A(net_7519), .ZN(net_642) );
SDFFR_X2 inst_2432 ( .D(net_4699), .SE(net_2313), .SI(net_404), .Q(net_404), .CK(net_16661), .RN(x6501) );
NAND2_X2 inst_4263 ( .A1(net_6913), .A2(net_5247), .ZN(net_5197) );
CLKBUF_X2 inst_14698 ( .A(net_14545), .Z(net_14546) );
HA_X1 inst_6693 ( .A(net_4459), .S(net_2873), .CO(net_2872), .B(net_2868) );
INV_X8 inst_5061 ( .ZN(net_6272), .A(net_4269) );
AOI22_X2 inst_8273 ( .B1(net_8728), .A1(net_8506), .ZN(net_6067), .B2(net_4350), .A2(net_4349) );
CLKBUF_X2 inst_10130 ( .A(net_9977), .Z(net_9978) );
NAND2_X2 inst_4343 ( .A1(net_7065), .A2(net_5162), .ZN(net_5114) );
AOI22_X2 inst_8560 ( .A1(net_2762), .B2(net_2556), .ZN(net_2456), .A2(net_2219), .B1(net_1936) );
CLKBUF_X2 inst_16352 ( .A(net_16199), .Z(net_16200) );
CLKBUF_X2 inst_15399 ( .A(net_15246), .Z(net_15247) );
INV_X4 inst_5684 ( .ZN(net_575), .A(net_275) );
CLKBUF_X2 inst_11537 ( .A(net_11384), .Z(net_11385) );
INV_X16 inst_6627 ( .ZN(net_4398), .A(net_3528) );
CLKBUF_X2 inst_11841 ( .A(net_10285), .Z(net_11689) );
XNOR2_X2 inst_235 ( .ZN(net_1245), .B(net_876), .A(net_517) );
CLKBUF_X2 inst_11493 ( .A(net_10146), .Z(net_11341) );
AOI222_X1 inst_8610 ( .B2(net_6769), .B1(net_5835), .A2(net_5830), .C2(net_5824), .ZN(net_5803), .A1(net_2822), .C1(net_2125) );
CLKBUF_X2 inst_12257 ( .A(net_12104), .Z(net_12105) );
INV_X4 inst_5643 ( .A(net_7615), .ZN(net_847) );
DFF_X1 inst_6750 ( .Q(net_6760), .D(net_5616), .CK(net_10497) );
CLKBUF_X2 inst_12555 ( .A(net_12170), .Z(net_12403) );
AOI22_X2 inst_8217 ( .B1(net_8758), .A1(net_8388), .A2(net_3867), .B2(net_3866), .ZN(net_3819) );
AOI22_X2 inst_8370 ( .B1(net_8744), .A1(net_8374), .A2(net_3867), .B2(net_3866), .ZN(net_3678) );
CLKBUF_X2 inst_12051 ( .A(net_11898), .Z(net_11899) );
NAND2_X2 inst_4338 ( .A1(net_7144), .A2(net_5166), .ZN(net_5119) );
AOI221_X2 inst_8806 ( .C2(net_5535), .B2(net_5260), .A(net_4898), .ZN(net_4722), .B1(net_3239), .C1(net_468) );
CLKBUF_X2 inst_16784 ( .A(net_16631), .Z(net_16632) );
AOI22_X2 inst_8194 ( .A1(net_8606), .B1(net_8421), .A2(net_3864), .B2(net_3863), .ZN(net_3841) );
OR2_X4 inst_2835 ( .A1(net_8901), .A2(net_6144), .ZN(net_4850) );
CLKBUF_X2 inst_12846 ( .A(net_12693), .Z(net_12694) );
CLKBUF_X2 inst_16907 ( .A(net_16754), .Z(net_16755) );
SDFFR_X1 inst_2731 ( .SI(net_9017), .Q(net_9017), .D(net_7446), .SE(net_3208), .CK(net_10109), .RN(x6501) );
CLKBUF_X2 inst_10399 ( .A(net_10246), .Z(net_10247) );
CLKBUF_X2 inst_11136 ( .A(net_10983), .Z(net_10984) );
AOI222_X1 inst_8663 ( .A2(net_3599), .B2(net_3598), .C2(net_3597), .ZN(net_3596), .A1(net_3595), .B1(net_1962), .C1(net_667) );
CLKBUF_X2 inst_17971 ( .A(net_9980), .Z(net_17819) );
NAND2_X2 inst_4813 ( .A2(net_2556), .ZN(net_1281), .A1(net_1280) );
CLKBUF_X2 inst_16960 ( .A(net_16807), .Z(net_16808) );
CLKBUF_X2 inst_9725 ( .A(net_9572), .Z(net_9573) );
CLKBUF_X2 inst_18488 ( .A(net_18335), .Z(net_18336) );
CLKBUF_X2 inst_15348 ( .A(net_15195), .Z(net_15196) );
CLKBUF_X2 inst_18178 ( .A(net_18025), .Z(net_18026) );
SDFF_X2 inst_477 ( .SI(net_8450), .Q(net_8450), .SE(net_3983), .D(net_3965), .CK(net_12466) );
NOR2_X2 inst_3398 ( .ZN(net_4562), .A1(net_4394), .A2(net_4368) );
NOR2_X2 inst_3576 ( .A1(net_5957), .ZN(net_1108), .A2(net_1106) );
SDFF_X2 inst_423 ( .SI(net_8306), .Q(net_8306), .SE(net_3978), .D(net_3946), .CK(net_11110) );
CLKBUF_X2 inst_10006 ( .A(net_9853), .Z(net_9854) );
CLKBUF_X2 inst_17367 ( .A(net_17214), .Z(net_17215) );
SDFF_X2 inst_835 ( .SI(net_8645), .Q(net_8645), .D(net_3973), .SE(net_3885), .CK(net_9981) );
OAI21_X2 inst_3082 ( .ZN(net_3156), .A(net_3154), .B2(net_3153), .B1(net_1167) );
NAND2_X2 inst_4137 ( .ZN(net_5384), .A1(net_5119), .A2(net_5118) );
DFF_X1 inst_6852 ( .Q(net_6440), .D(net_3628), .CK(net_17893) );
SDFF_X2 inst_1112 ( .D(net_7314), .SI(net_6523), .Q(net_6523), .SE(net_3086), .CK(net_9924) );
NAND2_X2 inst_4081 ( .A2(net_6786), .A1(net_5835), .ZN(net_5765) );
CLKBUF_X2 inst_9678 ( .A(net_9472), .Z(net_9526) );
CLKBUF_X2 inst_14571 ( .A(net_14418), .Z(net_14419) );
AOI21_X4 inst_8869 ( .B2(net_5948), .ZN(net_2486), .B1(net_2453), .A(net_2214) );
CLKBUF_X2 inst_18924 ( .A(net_18771), .Z(net_18772) );
SDFF_X2 inst_1817 ( .D(net_7294), .SI(net_6951), .Q(net_6951), .SE(net_6281), .CK(net_17683) );
CLKBUF_X2 inst_10375 ( .A(net_10222), .Z(net_10223) );
CLKBUF_X2 inst_17997 ( .A(net_17844), .Z(net_17845) );
CLKBUF_X2 inst_11056 ( .A(net_10903), .Z(net_10904) );
CLKBUF_X2 inst_19045 ( .A(net_18892), .Z(net_18893) );
CLKBUF_X2 inst_10081 ( .A(net_9928), .Z(net_9929) );
CLKBUF_X2 inst_14715 ( .A(net_14562), .Z(net_14563) );
OR2_X2 inst_2871 ( .A2(net_6132), .ZN(net_4780), .A1(net_1511) );
DFFR_X1 inst_7475 ( .QN(net_7431), .D(net_3992), .CK(net_12391), .RN(x6501) );
CLKBUF_X2 inst_17669 ( .A(net_17516), .Z(net_17517) );
NAND4_X2 inst_3629 ( .ZN(net_5583), .A1(net_5274), .A4(net_4810), .A3(net_4779), .A2(net_4477) );
CLKBUF_X2 inst_16297 ( .A(net_16144), .Z(net_16145) );
CLKBUF_X2 inst_12593 ( .A(net_12440), .Z(net_12441) );
CLKBUF_X2 inst_13370 ( .A(net_13217), .Z(net_13218) );
CLKBUF_X2 inst_9946 ( .A(net_9246), .Z(net_9794) );
CLKBUF_X2 inst_15427 ( .A(net_15274), .Z(net_15275) );
DFFR_X2 inst_7129 ( .QN(net_7600), .D(net_3084), .CK(net_9779), .RN(x6501) );
NAND2_X2 inst_4414 ( .A1(net_6853), .A2(net_5016), .ZN(net_5013) );
CLKBUF_X2 inst_18845 ( .A(net_18692), .Z(net_18693) );
CLKBUF_X2 inst_10052 ( .A(net_9899), .Z(net_9900) );
OAI21_X2 inst_3085 ( .ZN(net_3250), .B2(net_3033), .A(net_2951), .B1(net_1667) );
AOI222_X1 inst_8648 ( .A2(net_6266), .B2(net_4365), .C2(net_4364), .ZN(net_3918), .B1(net_3169), .C1(net_3167), .A1(x13722) );
CLKBUF_X2 inst_15337 ( .A(net_15184), .Z(net_15185) );
CLKBUF_X2 inst_16345 ( .A(net_16192), .Z(net_16193) );
CLKBUF_X2 inst_19005 ( .A(net_9183), .Z(net_18853) );
CLKBUF_X2 inst_16438 ( .A(net_10229), .Z(net_16286) );
CLKBUF_X2 inst_13768 ( .A(net_13615), .Z(net_13616) );
INV_X4 inst_5661 ( .A(net_7583), .ZN(net_581) );
CLKBUF_X2 inst_9918 ( .A(net_9065), .Z(net_9766) );
CLKBUF_X2 inst_11541 ( .A(net_11388), .Z(net_11389) );
CLKBUF_X2 inst_14120 ( .A(net_11424), .Z(net_13968) );
NAND2_X2 inst_4292 ( .A1(net_7040), .ZN(net_5168), .A2(net_5162) );
SDFFR_X2 inst_2449 ( .D(net_3111), .SE(net_2685), .SI(net_417), .Q(net_417), .CK(net_16894), .RN(x6501) );
CLKBUF_X2 inst_12083 ( .A(net_11757), .Z(net_11931) );
INV_X2 inst_6570 ( .A(net_6804), .ZN(net_487) );
CLKBUF_X2 inst_14709 ( .A(net_14556), .Z(net_14557) );
CLKBUF_X2 inst_13096 ( .A(net_10964), .Z(net_12944) );
SDFF_X2 inst_1431 ( .SI(net_7269), .Q(net_7046), .D(net_7046), .SE(net_6280), .CK(net_16860) );
NAND4_X2 inst_3760 ( .ZN(net_4261), .A1(net_3831), .A2(net_3830), .A3(net_3829), .A4(net_3828) );
SDFF_X2 inst_1398 ( .Q(net_8197), .D(net_8197), .SI(net_2719), .SE(net_2561), .CK(net_18802) );
CLKBUF_X2 inst_12841 ( .A(net_11498), .Z(net_12689) );
CLKBUF_X2 inst_18514 ( .A(net_17710), .Z(net_18362) );
DFFR_X2 inst_7122 ( .QN(net_7603), .D(net_3076), .CK(net_9789), .RN(x6501) );
AOI22_X2 inst_8477 ( .B1(net_6741), .A1(net_6708), .B2(net_6202), .A2(net_3520), .ZN(net_3463) );
OR2_X4 inst_2849 ( .A1(net_1910), .ZN(net_1739), .A2(net_1669) );
SDFFR_X2 inst_2440 ( .SE(net_2757), .D(net_2670), .SI(net_452), .Q(net_452), .CK(net_13829), .RN(x6501) );
CLKBUF_X2 inst_13808 ( .A(net_13655), .Z(net_13656) );
CLKBUF_X2 inst_9261 ( .A(net_9108), .Z(net_9109) );
CLKBUF_X2 inst_15533 ( .A(net_10700), .Z(net_15381) );
NOR2_X4 inst_3327 ( .ZN(net_3371), .A1(net_3260), .A2(net_3221) );
CLKBUF_X2 inst_10241 ( .A(net_10088), .Z(net_10089) );
SDFFR_X2 inst_2134 ( .SI(net_7202), .Q(net_7202), .D(net_6453), .SE(net_4362), .CK(net_16437), .RN(x6501) );
SDFF_X2 inst_1744 ( .Q(net_7905), .D(net_7905), .SI(net_2716), .SE(net_2543), .CK(net_16816) );
NAND2_X2 inst_4805 ( .ZN(net_1574), .A1(net_1334), .A2(net_1333) );
INV_X4 inst_5628 ( .A(net_7587), .ZN(net_588) );
CLKBUF_X2 inst_11958 ( .A(net_10561), .Z(net_11806) );
NAND2_X2 inst_4117 ( .ZN(net_5411), .A2(net_5232), .A1(net_5138) );
CLKBUF_X2 inst_11311 ( .A(net_11158), .Z(net_11159) );
CLKBUF_X2 inst_9329 ( .A(net_9176), .Z(net_9177) );
CLKBUF_X2 inst_10047 ( .A(net_9894), .Z(net_9895) );
CLKBUF_X2 inst_11198 ( .A(net_11045), .Z(net_11046) );
CLKBUF_X2 inst_11639 ( .A(net_10539), .Z(net_11487) );
CLKBUF_X2 inst_16480 ( .A(net_16327), .Z(net_16328) );
DFFS_X1 inst_6940 ( .D(net_6145), .CK(net_13646), .SN(x6501), .Q(x742) );
CLKBUF_X2 inst_11954 ( .A(net_9059), .Z(net_11802) );
CLKBUF_X2 inst_17354 ( .A(net_17201), .Z(net_17202) );
SDFF_X2 inst_712 ( .SI(net_8636), .Q(net_8636), .D(net_3947), .SE(net_3885), .CK(net_12961) );
CLKBUF_X2 inst_14271 ( .A(net_10496), .Z(net_14119) );
CLKBUF_X2 inst_12436 ( .A(net_12283), .Z(net_12284) );
OAI21_X2 inst_3111 ( .ZN(net_2477), .B2(net_2415), .B1(net_1860), .A(net_1586) );
CLKBUF_X2 inst_18455 ( .A(net_14518), .Z(net_18303) );
SDFF_X2 inst_2035 ( .SI(net_7915), .Q(net_7915), .D(net_2658), .SE(net_2461), .CK(net_15475) );
CLKBUF_X2 inst_17121 ( .A(net_10302), .Z(net_16969) );
CLKBUF_X2 inst_16500 ( .A(net_11508), .Z(net_16348) );
CLKBUF_X2 inst_13530 ( .A(net_13377), .Z(net_13378) );
CLKBUF_X2 inst_10442 ( .A(net_10289), .Z(net_10290) );
CLKBUF_X2 inst_11569 ( .A(net_10088), .Z(net_11417) );
CLKBUF_X2 inst_11121 ( .A(net_10968), .Z(net_10969) );
CLKBUF_X2 inst_14686 ( .A(net_12184), .Z(net_14534) );
CLKBUF_X2 inst_16252 ( .A(net_16099), .Z(net_16100) );
CLKBUF_X2 inst_17037 ( .A(net_16884), .Z(net_16885) );
CLKBUF_X2 inst_17023 ( .A(net_16870), .Z(net_16871) );
CLKBUF_X2 inst_12564 ( .A(net_12411), .Z(net_12412) );
CLKBUF_X2 inst_16782 ( .A(net_16137), .Z(net_16630) );
CLKBUF_X2 inst_16529 ( .A(net_11175), .Z(net_16377) );
INV_X2 inst_6483 ( .A(net_8269), .ZN(net_562) );
CLKBUF_X2 inst_12482 ( .A(net_12329), .Z(net_12330) );
DFFR_X1 inst_7381 ( .D(net_5894), .CK(net_11443), .RN(x6501), .Q(x2494) );
SDFF_X2 inst_525 ( .Q(net_8881), .D(net_8881), .SI(net_3952), .SE(net_3936), .CK(net_12900) );
CLKBUF_X2 inst_18735 ( .A(net_18582), .Z(net_18583) );
CLKBUF_X2 inst_17241 ( .A(net_13547), .Z(net_17089) );
CLKBUF_X2 inst_15360 ( .A(net_15207), .Z(net_15208) );
CLKBUF_X2 inst_11774 ( .A(net_11621), .Z(net_11622) );
CLKBUF_X2 inst_12196 ( .A(net_12043), .Z(net_12044) );
SDFF_X2 inst_1032 ( .SI(net_7317), .Q(net_6658), .D(net_6658), .SE(net_3126), .CK(net_12107) );
CLKBUF_X2 inst_12424 ( .A(net_12271), .Z(net_12272) );
AOI21_X2 inst_8985 ( .ZN(net_1889), .A(net_1888), .B2(net_1769), .B1(net_1454) );
HA_X1 inst_6711 ( .B(net_4360), .A(net_4355), .S(net_1235), .CO(net_1234) );
CLKBUF_X2 inst_12638 ( .A(net_11319), .Z(net_12486) );
CLKBUF_X2 inst_16580 ( .A(net_16427), .Z(net_16428) );
CLKBUF_X2 inst_18646 ( .A(net_18493), .Z(net_18494) );
INV_X4 inst_5932 ( .A(net_6289), .ZN(net_2675) );
CLKBUF_X2 inst_11682 ( .A(net_10925), .Z(net_11530) );
CLKBUF_X2 inst_11148 ( .A(net_10995), .Z(net_10996) );
CLKBUF_X2 inst_12339 ( .A(net_9887), .Z(net_12187) );
CLKBUF_X2 inst_11106 ( .A(net_10953), .Z(net_10954) );
CLKBUF_X2 inst_17413 ( .A(net_17260), .Z(net_17261) );
SDFFR_X2 inst_2269 ( .D(net_7385), .SE(net_2797), .SI(net_194), .Q(net_194), .CK(net_18153), .RN(x6501) );
SDFF_X2 inst_1780 ( .D(net_7280), .SI(net_6857), .Q(net_6857), .SE(net_6282), .CK(net_19017) );
CLKBUF_X2 inst_18459 ( .A(net_18306), .Z(net_18307) );
CLKBUF_X2 inst_11839 ( .A(net_11686), .Z(net_11687) );
SDFF_X2 inst_1436 ( .SI(net_7279), .Q(net_7096), .D(net_7096), .SE(net_6278), .CK(net_14638) );
SDFF_X2 inst_852 ( .SI(net_8665), .Q(net_8665), .D(net_3949), .SE(net_3885), .CK(net_12783) );
CLKBUF_X2 inst_12792 ( .A(net_11495), .Z(net_12640) );
HA_X1 inst_6663 ( .CO(net_6174), .S(net_3534), .A(net_3533), .B(net_3225) );
NAND2_X2 inst_4306 ( .A1(net_7094), .A2(net_5164), .ZN(net_5151) );
SDFF_X2 inst_1474 ( .SI(net_7268), .Q(net_7125), .D(net_7125), .SE(net_6279), .CK(net_17073) );
CLKBUF_X2 inst_12528 ( .A(net_12375), .Z(net_12376) );
CLKBUF_X2 inst_17821 ( .A(net_10807), .Z(net_17669) );
CLKBUF_X2 inst_11974 ( .A(net_11821), .Z(net_11822) );
CLKBUF_X2 inst_17563 ( .A(net_17410), .Z(net_17411) );
SDFF_X2 inst_1920 ( .D(net_7270), .SI(net_6847), .Q(net_6847), .SE(net_6282), .CK(net_14327) );
AOI211_X2 inst_9022 ( .C1(net_6111), .ZN(net_1429), .A(net_1324), .B(net_1322), .C2(net_1134) );
CLKBUF_X2 inst_19142 ( .A(net_18989), .Z(net_18990) );
CLKBUF_X2 inst_13269 ( .A(net_13116), .Z(net_13117) );
CLKBUF_X2 inst_18047 ( .A(net_17894), .Z(net_17895) );
CLKBUF_X2 inst_12787 ( .A(net_12411), .Z(net_12635) );
NAND2_X2 inst_4143 ( .ZN(net_5376), .A1(net_5113), .A2(net_5112) );
NOR4_X2 inst_3234 ( .ZN(net_1906), .A4(net_1651), .A2(net_1013), .A3(net_1009), .A1(net_965) );
CLKBUF_X2 inst_11194 ( .A(net_9541), .Z(net_11042) );
SDFFR_X2 inst_2639 ( .Q(net_7397), .D(net_2760), .SE(net_1136), .CK(net_14948), .RN(x6501), .SI(x4420) );
CLKBUF_X2 inst_18554 ( .A(net_12455), .Z(net_18402) );
CLKBUF_X2 inst_11122 ( .A(net_10969), .Z(net_10970) );
CLKBUF_X2 inst_15666 ( .A(net_10421), .Z(net_15514) );
INV_X4 inst_5897 ( .A(net_7231), .ZN(net_1855) );
INV_X16 inst_6632 ( .ZN(net_4349), .A(net_3368) );
SDFFR_X2 inst_2542 ( .QN(net_6368), .SE(net_2147), .SI(net_1867), .D(net_1241), .CK(net_18143), .RN(x6501) );
CLKBUF_X2 inst_15864 ( .A(net_15711), .Z(net_15712) );
CLKBUF_X2 inst_11791 ( .A(net_9293), .Z(net_11639) );
DFF_X1 inst_6829 ( .Q(net_6449), .D(net_3619), .CK(net_17912) );
CLKBUF_X2 inst_9506 ( .A(net_9353), .Z(net_9354) );
DFFR_X1 inst_7567 ( .Q(net_6825), .D(net_6813), .CK(net_15125), .RN(x6501) );
INV_X2 inst_6590 ( .A(net_6120), .ZN(net_6119) );
SDFF_X2 inst_417 ( .SI(net_8332), .Q(net_8332), .SE(net_3978), .D(net_3949), .CK(net_10589) );
SDFF_X2 inst_671 ( .Q(net_8415), .D(net_8415), .SI(net_3981), .SE(net_3934), .CK(net_12966) );
CLKBUF_X2 inst_18356 ( .A(net_18203), .Z(net_18204) );
CLKBUF_X2 inst_12733 ( .A(net_12580), .Z(net_12581) );
CLKBUF_X2 inst_13473 ( .A(net_13320), .Z(net_13321) );
CLKBUF_X2 inst_15812 ( .A(net_15659), .Z(net_15660) );
CLKBUF_X2 inst_18083 ( .A(net_17001), .Z(net_17931) );
XOR2_X2 inst_21 ( .Z(net_1398), .B(net_1397), .A(net_647) );
CLKBUF_X2 inst_9462 ( .A(net_9113), .Z(net_9310) );
CLKBUF_X2 inst_14782 ( .A(net_14629), .Z(net_14630) );
CLKBUF_X2 inst_18364 ( .A(net_11264), .Z(net_18212) );
CLKBUF_X2 inst_17724 ( .A(net_13056), .Z(net_17572) );
CLKBUF_X2 inst_18741 ( .A(net_15052), .Z(net_18589) );
CLKBUF_X2 inst_16381 ( .A(net_16228), .Z(net_16229) );
CLKBUF_X2 inst_11024 ( .A(net_9092), .Z(net_10872) );
CLKBUF_X2 inst_10286 ( .A(net_10133), .Z(net_10134) );
CLKBUF_X2 inst_19163 ( .A(net_19010), .Z(net_19011) );
SDFFR_X2 inst_2311 ( .SE(net_2260), .Q(net_378), .D(net_378), .CK(net_11475), .RN(x6501), .SI(x1383) );
NAND3_X2 inst_3885 ( .ZN(net_5886), .A3(net_5773), .A1(net_4960), .A2(net_4781) );
CLKBUF_X2 inst_17309 ( .A(net_13096), .Z(net_17157) );
NAND4_X2 inst_3683 ( .A4(net_6240), .A1(net_6239), .ZN(net_4454), .A2(net_3873), .A3(net_3872) );
OAI22_X2 inst_2941 ( .A1(net_2097), .ZN(net_1879), .B1(net_1778), .A2(net_1616), .B2(net_1327) );
CLKBUF_X2 inst_13655 ( .A(net_13502), .Z(net_13503) );
CLKBUF_X2 inst_13528 ( .A(net_13375), .Z(net_13376) );
CLKBUF_X2 inst_9861 ( .A(net_9324), .Z(net_9709) );
CLKBUF_X2 inst_12351 ( .A(net_12198), .Z(net_12199) );
AND2_X2 inst_9203 ( .ZN(net_6062), .A1(net_904), .A2(net_903) );
AOI22_X2 inst_8442 ( .B1(net_6733), .A1(net_6700), .B2(net_6202), .A2(net_3520), .ZN(net_3499) );
CLKBUF_X2 inst_17742 ( .A(net_17589), .Z(net_17590) );
CLKBUF_X2 inst_10920 ( .A(net_10303), .Z(net_10768) );
CLKBUF_X2 inst_11930 ( .A(net_11777), .Z(net_11778) );
CLKBUF_X2 inst_18618 ( .A(net_11243), .Z(net_18466) );
SDFFR_X2 inst_2637 ( .Q(net_7372), .D(net_7372), .SE(net_1136), .CK(net_18601), .RN(x6501), .SI(x4805) );
CLKBUF_X2 inst_9604 ( .A(net_9451), .Z(net_9452) );
CLKBUF_X2 inst_16319 ( .A(net_16166), .Z(net_16167) );
XNOR2_X2 inst_236 ( .ZN(net_1242), .A(net_1241), .B(net_879) );
NAND2_X2 inst_4539 ( .A1(net_3374), .ZN(net_3368), .A2(net_3367) );
NAND3_X4 inst_3878 ( .ZN(net_2027), .A3(net_1562), .A2(net_1530), .A1(net_1498) );
CLKBUF_X2 inst_13295 ( .A(net_13142), .Z(net_13143) );
CLKBUF_X2 inst_9806 ( .A(net_9653), .Z(net_9654) );
SDFF_X2 inst_986 ( .D(net_7323), .SI(net_6631), .Q(net_6631), .SE(net_3123), .CK(net_11357) );
OAI21_X2 inst_3172 ( .B1(net_9004), .A(net_1886), .ZN(net_1059), .B2(net_767) );
MUX2_X2 inst_4983 ( .A(net_9032), .Z(net_3967), .B(net_3170), .S(net_622) );
SDFF_X2 inst_1422 ( .SI(net_7278), .Q(net_7055), .D(net_7055), .SE(net_6280), .CK(net_14643) );
CLKBUF_X2 inst_10263 ( .A(net_9927), .Z(net_10111) );
AOI22_X2 inst_8337 ( .B1(net_8773), .A1(net_8403), .A2(net_3867), .B2(net_3866), .ZN(net_3710) );
CLKBUF_X2 inst_9702 ( .A(net_9075), .Z(net_9550) );
DFFS_X2 inst_6893 ( .QN(net_8969), .D(net_2856), .CK(net_17612), .SN(x6501) );
CLKBUF_X2 inst_10522 ( .A(net_10369), .Z(net_10370) );
SDFF_X2 inst_1221 ( .Q(net_7952), .D(net_7952), .SE(net_2755), .SI(net_2584), .CK(net_16089) );
AOI222_X1 inst_8675 ( .C2(net_5832), .A2(net_5830), .B2(net_5824), .ZN(net_3361), .A1(net_3166), .B1(net_2120), .C1(x2400) );
CLKBUF_X2 inst_19149 ( .A(net_15598), .Z(net_18997) );
AOI22_X2 inst_7750 ( .B1(net_6979), .A1(net_6939), .A2(net_5443), .B2(net_5442), .ZN(net_5406) );
CLKBUF_X2 inst_12158 ( .A(net_12005), .Z(net_12006) );
CLKBUF_X2 inst_15000 ( .A(net_14847), .Z(net_14848) );
AOI22_X2 inst_7951 ( .B1(net_8192), .A1(net_7682), .B2(net_6099), .A2(net_4399), .ZN(net_4175) );
CLKBUF_X2 inst_16005 ( .A(net_14587), .Z(net_15853) );
CLKBUF_X2 inst_15121 ( .A(net_14968), .Z(net_14969) );
INV_X4 inst_5139 ( .ZN(net_3557), .A(net_3527) );
CLKBUF_X2 inst_16240 ( .A(net_16087), .Z(net_16088) );
SDFFR_X1 inst_2664 ( .D(net_6761), .SE(net_4506), .CK(net_11539), .RN(x6501), .SI(x2041), .Q(x2041) );
CLKBUF_X2 inst_10793 ( .A(net_10640), .Z(net_10641) );
AOI221_X2 inst_8761 ( .C2(net_6130), .B2(net_5535), .ZN(net_5471), .A(net_4947), .C1(net_1387), .B1(net_461) );
CLKBUF_X2 inst_11615 ( .A(net_11462), .Z(net_11463) );
CLKBUF_X2 inst_15463 ( .A(net_15310), .Z(net_15311) );
DFF_X1 inst_6757 ( .Q(net_7537), .D(net_4615), .CK(net_11981) );
CLKBUF_X2 inst_19197 ( .A(net_12194), .Z(net_19045) );
AOI22_X2 inst_8170 ( .B1(net_8788), .A1(net_8529), .ZN(net_3862), .A2(net_3861), .B2(net_3860) );
AOI22_X2 inst_7915 ( .A2(net_6427), .A1(net_5654), .ZN(net_4488), .B2(net_4486), .B1(net_264) );
INV_X4 inst_5862 ( .A(net_6309), .ZN(net_2681) );
CLKBUF_X2 inst_14007 ( .A(net_12700), .Z(net_13855) );
CLKBUF_X2 inst_19138 ( .A(net_13168), .Z(net_18986) );
CLKBUF_X2 inst_10966 ( .A(net_10813), .Z(net_10814) );
CLKBUF_X2 inst_18080 ( .A(net_17927), .Z(net_17928) );
CLKBUF_X2 inst_11381 ( .A(net_11228), .Z(net_11229) );
CLKBUF_X2 inst_15253 ( .A(net_14143), .Z(net_15101) );
CLKBUF_X2 inst_10570 ( .A(net_10417), .Z(net_10418) );
AOI22_X2 inst_8051 ( .B1(net_8206), .A1(net_7696), .B2(net_6099), .A2(net_4399), .ZN(net_4090) );
AOI22_X2 inst_8413 ( .B1(net_8787), .A1(net_8528), .A2(net_3861), .B2(net_3860), .ZN(net_3639) );
CLKBUF_X2 inst_16090 ( .A(net_15937), .Z(net_15938) );
NAND3_X2 inst_3932 ( .ZN(net_5529), .A1(net_5262), .A3(net_4733), .A2(net_4651) );
CLKBUF_X2 inst_15811 ( .A(net_15658), .Z(net_15659) );
CLKBUF_X2 inst_16162 ( .A(net_13722), .Z(net_16010) );
CLKBUF_X2 inst_16520 ( .A(net_13155), .Z(net_16368) );
CLKBUF_X2 inst_13634 ( .A(net_13481), .Z(net_13482) );
INV_X2 inst_6295 ( .ZN(net_4203), .A(net_3912) );
CLKBUF_X2 inst_16736 ( .A(net_9871), .Z(net_16584) );
CLKBUF_X2 inst_17323 ( .A(net_17170), .Z(net_17171) );
CLKBUF_X2 inst_11433 ( .A(net_10666), .Z(net_11281) );
CLKBUF_X2 inst_11429 ( .A(net_11276), .Z(net_11277) );
CLKBUF_X2 inst_18136 ( .A(net_17983), .Z(net_17984) );
CLKBUF_X2 inst_18590 ( .A(net_18437), .Z(net_18438) );
CLKBUF_X2 inst_15980 ( .A(net_15827), .Z(net_15828) );
INV_X4 inst_5512 ( .ZN(net_682), .A(net_681) );
CLKBUF_X2 inst_13112 ( .A(net_12959), .Z(net_12960) );
CLKBUF_X2 inst_11973 ( .A(net_11820), .Z(net_11821) );
CLKBUF_X2 inst_12265 ( .A(net_9329), .Z(net_12113) );
NAND4_X2 inst_3781 ( .ZN(net_4240), .A1(net_3698), .A2(net_3697), .A3(net_3696), .A4(net_3695) );
AND2_X4 inst_9081 ( .ZN(net_3126), .A2(net_2940), .A1(net_2902) );
NOR2_X2 inst_3552 ( .ZN(net_2071), .A1(net_1591), .A2(net_1475) );
SDFF_X2 inst_1702 ( .Q(net_8205), .D(net_8205), .SI(net_2711), .SE(net_2561), .CK(net_14162) );
SDFF_X2 inst_1277 ( .Q(net_8110), .D(net_8110), .SE(net_2707), .SI(net_2656), .CK(net_14028) );
CLKBUF_X2 inst_17802 ( .A(net_17649), .Z(net_17650) );
NAND2_X2 inst_4076 ( .A2(net_6774), .A1(net_5835), .ZN(net_5770) );
SDFFS_X2 inst_2092 ( .SI(net_6828), .Q(net_6828), .SE(net_2146), .D(net_2104), .CK(net_18672), .SN(x6501) );
INV_X4 inst_5586 ( .A(net_6469), .ZN(net_1202) );
CLKBUF_X2 inst_13784 ( .A(net_13631), .Z(net_13632) );
SDFF_X2 inst_1440 ( .SI(net_7283), .Q(net_7100), .D(net_7100), .SE(net_6278), .CK(net_16225) );
CLKBUF_X2 inst_9415 ( .A(net_9238), .Z(net_9263) );
CLKBUF_X2 inst_13611 ( .A(net_12676), .Z(net_13459) );
CLKBUF_X2 inst_15522 ( .A(net_15369), .Z(net_15370) );
CLKBUF_X2 inst_9854 ( .A(net_9701), .Z(net_9702) );
CLKBUF_X2 inst_13734 ( .A(net_13581), .Z(net_13582) );
NOR2_X2 inst_3355 ( .ZN(net_5570), .A1(net_5408), .A2(net_5407) );
CLKBUF_X2 inst_12148 ( .A(net_10535), .Z(net_11996) );
AOI22_X2 inst_8179 ( .B1(net_8826), .A1(net_8345), .A2(net_6265), .B2(net_6253), .ZN(net_6076) );
INV_X2 inst_6213 ( .ZN(net_5497), .A(net_5377) );
CLKBUF_X2 inst_17214 ( .A(net_17061), .Z(net_17062) );
AOI22_X2 inst_8354 ( .B1(net_8850), .A1(net_8369), .A2(net_6265), .B2(net_6253), .ZN(net_3694) );
SDFF_X2 inst_1591 ( .Q(net_8122), .D(net_8122), .SI(net_2584), .SE(net_2541), .CK(net_18380) );
NAND4_X2 inst_3697 ( .ZN(net_4440), .A4(net_4341), .A1(net_3782), .A2(net_3781), .A3(net_3780) );
INV_X4 inst_5470 ( .ZN(net_752), .A(net_751) );
AOI22_X2 inst_7827 ( .A2(net_5657), .B2(net_5535), .ZN(net_4694), .A1(net_2695), .B1(net_450) );
AOI22_X2 inst_8312 ( .B1(net_8817), .A1(net_8336), .A2(net_6265), .B2(net_6253), .ZN(net_3733) );
SDFFR_X2 inst_2570 ( .QN(net_6376), .SE(net_2147), .D(net_2120), .SI(net_1958), .CK(net_18128), .RN(x6501) );
CLKBUF_X2 inst_12856 ( .A(net_12703), .Z(net_12704) );
CLKBUF_X2 inst_18375 ( .A(net_18222), .Z(net_18223) );
MUX2_X2 inst_4960 ( .A(net_7379), .S(net_2376), .Z(net_2363), .B(net_800) );
CLKBUF_X2 inst_16811 ( .A(net_16658), .Z(net_16659) );
CLKBUF_X2 inst_14205 ( .A(net_14052), .Z(net_14053) );
AND2_X4 inst_9098 ( .ZN(net_2545), .A2(net_2268), .A1(net_2263) );
NAND4_X2 inst_3719 ( .ZN(net_4418), .A4(net_4327), .A1(net_3642), .A2(net_3641), .A3(net_3640) );
NAND2_X2 inst_4095 ( .ZN(net_5440), .A1(net_5161), .A2(net_5160) );
XOR2_X1 inst_74 ( .Z(net_3331), .B(net_3330), .A(net_3195) );
CLKBUF_X2 inst_15926 ( .A(net_13516), .Z(net_15774) );
SDFFR_X2 inst_2244 ( .SE(net_2814), .SI(net_2803), .Q(net_245), .D(net_245), .CK(net_14718), .RN(x6501) );
CLKBUF_X2 inst_13357 ( .A(net_12643), .Z(net_13205) );
CLKBUF_X2 inst_18760 ( .A(net_18607), .Z(net_18608) );
CLKBUF_X2 inst_14739 ( .A(net_11520), .Z(net_14587) );
NOR3_X2 inst_3284 ( .ZN(net_2732), .A1(net_2400), .A3(net_2319), .A2(net_1140) );
CLKBUF_X2 inst_11435 ( .A(net_11282), .Z(net_11283) );
CLKBUF_X2 inst_18652 ( .A(net_18499), .Z(net_18500) );
INV_X4 inst_5719 ( .A(net_8936), .ZN(net_2600) );
INV_X4 inst_5648 ( .A(net_7569), .ZN(net_586) );
NAND2_X2 inst_4512 ( .A2(net_6212), .ZN(net_4370), .A1(net_4274) );
CLKBUF_X2 inst_14265 ( .A(net_14112), .Z(net_14113) );
CLKBUF_X2 inst_16946 ( .A(net_16793), .Z(net_16794) );
AOI22_X2 inst_8483 ( .B1(net_6610), .A1(net_6577), .A2(net_6257), .B2(net_6110), .ZN(net_3457) );
CLKBUF_X2 inst_18936 ( .A(net_18783), .Z(net_18784) );
INV_X4 inst_5991 ( .A(net_5969), .ZN(x3258) );
CLKBUF_X2 inst_11234 ( .A(net_11081), .Z(net_11082) );
CLKBUF_X2 inst_13619 ( .A(net_10670), .Z(net_13467) );
DFFS_X1 inst_6949 ( .D(net_6145), .CK(net_16342), .SN(x6501), .Q(x838) );
CLKBUF_X2 inst_17919 ( .A(net_17766), .Z(net_17767) );
CLKBUF_X2 inst_16506 ( .A(net_14810), .Z(net_16354) );
INV_X4 inst_5709 ( .ZN(net_762), .A(net_401) );
CLKBUF_X2 inst_11401 ( .A(net_11248), .Z(net_11249) );
CLKBUF_X2 inst_16573 ( .A(net_11469), .Z(net_16421) );
INV_X4 inst_5335 ( .ZN(net_1454), .A(net_1335) );
SDFFR_X2 inst_2397 ( .SI(net_2785), .SE(net_2723), .D(net_2699), .QN(net_162), .CK(net_15038), .RN(x6501) );
CLKBUF_X2 inst_12802 ( .A(net_12649), .Z(net_12650) );
CLKBUF_X2 inst_13539 ( .A(net_9507), .Z(net_13387) );
SDFF_X2 inst_1090 ( .D(net_7315), .SI(net_6491), .Q(net_6491), .SE(net_3071), .CK(net_12089) );
CLKBUF_X2 inst_9709 ( .A(net_9556), .Z(net_9557) );
AND2_X4 inst_9088 ( .A1(net_2741), .ZN(net_2582), .A2(net_2475) );
SDFFR_X2 inst_2372 ( .SE(net_2260), .Q(net_307), .D(net_307), .CK(net_9297), .RN(x6501), .SI(x3651) );
SDFFR_X2 inst_2575 ( .D(net_7383), .QN(net_7243), .SI(net_1961), .SE(net_1379), .CK(net_18121), .RN(x6501) );
CLKBUF_X2 inst_17437 ( .A(net_9456), .Z(net_17285) );
MUX2_X2 inst_5007 ( .B(net_6324), .Z(net_4924), .S(net_644), .A(x4964) );
CLKBUF_X2 inst_10923 ( .A(net_10723), .Z(net_10771) );
CLKBUF_X2 inst_12496 ( .A(net_12343), .Z(net_12344) );
CLKBUF_X2 inst_13521 ( .A(net_13368), .Z(net_13369) );
INV_X4 inst_5655 ( .A(net_6820), .ZN(net_1216) );
CLKBUF_X2 inst_17071 ( .A(net_16918), .Z(net_16919) );
CLKBUF_X2 inst_16534 ( .A(net_10739), .Z(net_16382) );
CLKBUF_X2 inst_11874 ( .A(net_11721), .Z(net_11722) );
INV_X4 inst_5874 ( .A(net_8915), .ZN(net_2618) );
OAI21_X2 inst_3126 ( .A(net_2304), .ZN(net_2219), .B2(net_2122), .B1(net_1937) );
CLKBUF_X2 inst_12547 ( .A(net_12394), .Z(net_12395) );
AOI22_X2 inst_8028 ( .B1(net_8202), .A1(net_7692), .B2(net_6099), .A2(net_4399), .ZN(net_4109) );
SDFF_X2 inst_503 ( .SI(net_8596), .Q(net_8596), .SE(net_3984), .D(net_3977), .CK(net_10767) );
AOI221_X2 inst_8770 ( .C1(net_8986), .B2(net_5538), .C2(net_5456), .ZN(net_5278), .A(net_4874), .B1(net_415) );
CLKBUF_X2 inst_12107 ( .A(net_11954), .Z(net_11955) );
INV_X4 inst_5340 ( .ZN(net_4323), .A(net_1369) );
AOI221_X4 inst_8724 ( .B1(net_8837), .C1(net_8356), .C2(net_6265), .B2(net_6253), .ZN(net_4341), .A(net_4253) );
SDFF_X2 inst_1936 ( .SI(net_8067), .Q(net_8067), .D(net_2749), .SE(net_2508), .CK(net_16458) );
OAI211_X2 inst_3193 ( .ZN(net_3188), .A(net_3163), .B(net_3162), .C2(net_2067), .C1(net_1502) );
INV_X2 inst_6458 ( .A(net_8951), .ZN(net_790) );
SDFFS_X1 inst_2099 ( .SI(net_6810), .Q(net_6810), .SE(net_6267), .D(net_4622), .CK(net_11776), .SN(x6501) );
NAND2_X2 inst_4069 ( .A1(net_6335), .A2(net_6331), .ZN(net_5920) );
INV_X4 inst_5433 ( .A(net_863), .ZN(net_830) );
SDFF_X2 inst_1097 ( .D(net_7324), .SI(net_6533), .Q(net_6533), .SE(net_3086), .CK(net_9843) );
CLKBUF_X2 inst_11079 ( .A(net_9675), .Z(net_10927) );
CLKBUF_X2 inst_15268 ( .A(net_14203), .Z(net_15116) );
CLKBUF_X2 inst_16710 ( .A(net_16557), .Z(net_16558) );
OR2_X2 inst_2888 ( .ZN(net_1709), .A1(net_1685), .A2(net_1379) );
DFF_X1 inst_6804 ( .Q(net_8221), .D(net_4424), .CK(net_16565) );
CLKBUF_X2 inst_9382 ( .A(net_9069), .Z(net_9230) );
CLKBUF_X2 inst_12633 ( .A(net_9321), .Z(net_12481) );
CLKBUF_X2 inst_12683 ( .A(net_12530), .Z(net_12531) );
CLKBUF_X2 inst_12330 ( .A(net_12177), .Z(net_12178) );
SDFF_X2 inst_967 ( .SI(net_7328), .Q(net_6735), .D(net_6735), .SE(net_3124), .CK(net_9529) );
CLKBUF_X2 inst_9235 ( .A(net_9082), .Z(net_9083) );
CLKBUF_X2 inst_13117 ( .A(net_12964), .Z(net_12965) );
CLKBUF_X2 inst_18619 ( .A(net_10011), .Z(net_18467) );
CLKBUF_X2 inst_12665 ( .A(net_12512), .Z(net_12513) );
CLKBUF_X2 inst_16553 ( .A(net_16400), .Z(net_16401) );
AOI22_X2 inst_7863 ( .B2(net_5609), .A2(net_5267), .ZN(net_4578), .B1(net_376), .A1(net_180) );
CLKBUF_X2 inst_11495 ( .A(net_11342), .Z(net_11343) );
CLKBUF_X2 inst_12200 ( .A(net_12047), .Z(net_12048) );
CLKBUF_X2 inst_12029 ( .A(net_11876), .Z(net_11877) );
SDFF_X2 inst_1227 ( .Q(net_7958), .D(net_7958), .SE(net_2755), .SI(net_2575), .CK(net_16011) );
CLKBUF_X2 inst_16469 ( .A(net_16316), .Z(net_16317) );
CLKBUF_X2 inst_16522 ( .A(net_16369), .Z(net_16370) );
SDFFR_X2 inst_2324 ( .SE(net_2260), .Q(net_377), .D(net_377), .CK(net_11397), .RN(x6501), .SI(x1428) );
INV_X4 inst_5856 ( .A(net_7214), .ZN(net_1622) );
CLKBUF_X2 inst_9443 ( .A(net_9290), .Z(net_9291) );
INV_X4 inst_5732 ( .A(net_7239), .ZN(net_1941) );
OR2_X2 inst_2897 ( .A2(net_9053), .ZN(net_5990), .A1(net_895) );
CLKBUF_X2 inst_15086 ( .A(net_14676), .Z(net_14934) );
SDFFR_X2 inst_2529 ( .Q(net_7667), .D(net_7667), .SE(net_2299), .SI(net_1964), .CK(net_17262), .RN(x6501) );
CLKBUF_X2 inst_15687 ( .A(net_15534), .Z(net_15535) );
CLKBUF_X2 inst_11807 ( .A(net_11153), .Z(net_11655) );
SDFF_X2 inst_1787 ( .D(net_7282), .SI(net_6939), .Q(net_6939), .SE(net_6281), .CK(net_16203) );
CLKBUF_X2 inst_19087 ( .A(net_18934), .Z(net_18935) );
DFFR_X2 inst_7274 ( .QN(net_7357), .D(net_1901), .CK(net_11609), .RN(x6501) );
CLKBUF_X2 inst_12581 ( .A(net_12428), .Z(net_12429) );
CLKBUF_X2 inst_9741 ( .A(net_9380), .Z(net_9589) );
CLKBUF_X2 inst_14290 ( .A(net_9177), .Z(net_14138) );
INV_X4 inst_5943 ( .A(net_7495), .ZN(net_2916) );
CLKBUF_X2 inst_17844 ( .A(net_17691), .Z(net_17692) );
CLKBUF_X2 inst_9891 ( .A(net_9738), .Z(net_9739) );
INV_X2 inst_6310 ( .ZN(net_3894), .A(net_3591) );
SDFF_X2 inst_1540 ( .Q(net_7994), .D(net_7994), .SI(net_2590), .SE(net_2542), .CK(net_15591) );
CLKBUF_X2 inst_9493 ( .A(net_9089), .Z(net_9341) );
SDFFR_X1 inst_2742 ( .SI(net_9018), .Q(net_9018), .D(net_7447), .SE(net_3208), .CK(net_12836), .RN(x6501) );
NOR2_X2 inst_3536 ( .ZN(net_1571), .A2(net_1565), .A1(x13208) );
DFFR_X1 inst_7515 ( .Q(net_7310), .D(net_1664), .CK(net_9675), .RN(x6501) );
INV_X4 inst_5243 ( .ZN(net_2849), .A(net_1913) );
CLKBUF_X2 inst_12355 ( .A(net_9211), .Z(net_12203) );
SDFFR_X2 inst_2346 ( .SE(net_2260), .Q(net_310), .D(net_310), .CK(net_10466), .RN(x6501), .SI(x3524) );
CLKBUF_X2 inst_12486 ( .A(net_12333), .Z(net_12334) );
CLKBUF_X2 inst_12123 ( .A(net_11970), .Z(net_11971) );
CLKBUF_X2 inst_13653 ( .A(net_12238), .Z(net_13501) );
CLKBUF_X2 inst_15629 ( .A(net_15476), .Z(net_15477) );
DFFR_X2 inst_7250 ( .QN(net_7226), .D(net_2064), .CK(net_15048), .RN(x6501) );
CLKBUF_X2 inst_12291 ( .A(net_12138), .Z(net_12139) );
CLKBUF_X2 inst_15680 ( .A(net_10724), .Z(net_15528) );
DFFR_X2 inst_7363 ( .Q(net_7322), .CK(net_11757), .D(x13077), .RN(x6501) );
CLKBUF_X2 inst_9746 ( .A(net_9593), .Z(net_9594) );
CLKBUF_X2 inst_15279 ( .A(net_15126), .Z(net_15127) );
CLKBUF_X2 inst_17492 ( .A(net_17339), .Z(net_17340) );
CLKBUF_X2 inst_15135 ( .A(net_9136), .Z(net_14983) );
CLKBUF_X2 inst_16801 ( .A(net_16648), .Z(net_16649) );
DFFR_X2 inst_7171 ( .QN(net_7363), .D(net_2743), .CK(net_9510), .RN(x6501) );
SDFF_X2 inst_1005 ( .D(net_7316), .SI(net_6624), .Q(net_6624), .SE(net_3123), .CK(net_9872) );
CLKBUF_X2 inst_18767 ( .A(net_18614), .Z(net_18615) );
DFFR_X2 inst_6979 ( .QN(net_6293), .D(net_5914), .CK(net_16758), .RN(x6501) );
CLKBUF_X2 inst_14895 ( .A(net_14742), .Z(net_14743) );
SDFF_X2 inst_1580 ( .Q(net_8032), .D(net_8032), .SI(net_2712), .SE(net_2545), .CK(net_17139) );
SDFF_X2 inst_1842 ( .D(net_7278), .SI(net_6855), .Q(net_6855), .SE(net_6282), .CK(net_18996) );
CLKBUF_X2 inst_17456 ( .A(net_17303), .Z(net_17304) );
CLKBUF_X2 inst_17929 ( .A(net_14259), .Z(net_17777) );
DFFR_X1 inst_7534 ( .D(net_2695), .Q(net_294), .CK(net_11638), .RN(x6501) );
DFF_X1 inst_6737 ( .Q(net_6782), .D(net_5632), .CK(net_11428) );
NAND4_X2 inst_3703 ( .A4(net_6230), .A1(net_6229), .ZN(net_4434), .A2(net_3744), .A3(net_3743) );
SDFF_X2 inst_1333 ( .SI(net_7682), .Q(net_7682), .SE(net_2714), .D(net_2574), .CK(net_15619) );
CLKBUF_X2 inst_12613 ( .A(net_10769), .Z(net_12461) );
NAND3_X2 inst_3953 ( .A3(net_3533), .A2(net_3224), .ZN(net_3193), .A1(net_3192) );
DFFR_X2 inst_7315 ( .QN(net_6467), .D(net_6464), .CK(net_15096), .RN(x6501) );
SDFF_X2 inst_1551 ( .Q(net_8008), .D(net_8008), .SI(net_2656), .SE(net_2542), .CK(net_16720) );
CLKBUF_X2 inst_14505 ( .A(net_12191), .Z(net_14353) );
CLKBUF_X2 inst_9579 ( .A(net_9378), .Z(net_9427) );
SDFF_X2 inst_1088 ( .D(net_7342), .SI(net_6518), .Q(net_6518), .SE(net_3071), .CK(net_11678) );
CLKBUF_X2 inst_13200 ( .A(net_13047), .Z(net_13048) );
CLKBUF_X2 inst_15238 ( .A(net_15085), .Z(net_15086) );
AOI222_X1 inst_8692 ( .C2(net_5832), .A2(net_5830), .B2(net_5824), .ZN(net_3234), .A1(net_3091), .B1(net_2136), .C1(x3207) );
CLKBUF_X2 inst_15498 ( .A(net_15345), .Z(net_15346) );
CLKBUF_X2 inst_11672 ( .A(net_9606), .Z(net_11520) );
CLKBUF_X2 inst_13165 ( .A(net_13012), .Z(net_13013) );
INV_X4 inst_5844 ( .A(net_7387), .ZN(net_927) );
AOI221_X2 inst_8781 ( .B1(net_7188), .C2(net_6187), .B2(net_5655), .ZN(net_5257), .A(net_4933), .C1(net_189) );
CLKBUF_X2 inst_13142 ( .A(net_11471), .Z(net_12990) );
INV_X2 inst_6433 ( .ZN(net_691), .A(net_690) );
CLKBUF_X2 inst_9922 ( .A(net_9739), .Z(net_9770) );
CLKBUF_X2 inst_12941 ( .A(net_12788), .Z(net_12789) );
OAI22_X2 inst_2931 ( .B1(net_7225), .ZN(net_2448), .A2(net_2447), .B2(net_2063), .A1(net_1871) );
CLKBUF_X2 inst_18795 ( .A(net_18642), .Z(net_18643) );
NAND2_X2 inst_4768 ( .ZN(net_1766), .A2(net_1678), .A1(net_570) );
CLKBUF_X2 inst_14483 ( .A(net_14330), .Z(net_14331) );
SDFFR_X2 inst_2530 ( .Q(net_6412), .D(net_6412), .SI(net_6411), .SE(net_1893), .CK(net_17943), .RN(x6501) );
SDFF_X2 inst_1503 ( .SI(net_7862), .Q(net_7862), .D(net_2712), .SE(net_2558), .CK(net_13778) );
CLKBUF_X2 inst_12234 ( .A(net_12081), .Z(net_12082) );
INV_X4 inst_5656 ( .ZN(net_583), .A(net_270) );
AOI22_X2 inst_7874 ( .A2(net_6439), .A1(net_5654), .B2(net_4881), .ZN(net_4567), .B1(net_239) );
NAND4_X2 inst_3802 ( .ZN(net_3624), .A1(net_3479), .A2(net_3478), .A4(net_3477), .A3(net_3476) );
AOI22_X2 inst_8317 ( .B1(net_8669), .A1(net_8632), .B2(net_6109), .A2(net_3857), .ZN(net_3728) );
CLKBUF_X2 inst_12926 ( .A(net_9234), .Z(net_12774) );
CLKBUF_X2 inst_10718 ( .A(net_10565), .Z(net_10566) );
CLKBUF_X2 inst_11094 ( .A(net_10467), .Z(net_10942) );
SDFF_X2 inst_933 ( .SI(net_7313), .Q(net_6654), .D(net_6654), .SE(net_3126), .CK(net_12055) );
CLKBUF_X2 inst_13902 ( .A(net_13027), .Z(net_13750) );
CLKBUF_X2 inst_17566 ( .A(net_14202), .Z(net_17414) );
SDFF_X2 inst_1013 ( .SI(net_7327), .Q(net_6668), .D(net_6668), .SE(net_3126), .CK(net_9100) );
CLKBUF_X2 inst_14362 ( .A(net_14209), .Z(net_14210) );
NOR2_X2 inst_3613 ( .A2(net_7526), .A1(net_7522), .ZN(net_1430) );
CLKBUF_X2 inst_9439 ( .A(net_9286), .Z(net_9287) );
AOI22_X2 inst_7790 ( .A2(net_6187), .ZN(net_4810), .B2(net_4809), .B1(net_345), .A1(net_201) );
CLKBUF_X2 inst_12870 ( .A(net_12717), .Z(net_12718) );
CLKBUF_X2 inst_14054 ( .A(net_13901), .Z(net_13902) );
AOI22_X2 inst_8481 ( .B1(net_6742), .A1(net_6709), .B2(net_6202), .A2(net_3520), .ZN(net_3459) );
XNOR2_X2 inst_124 ( .ZN(net_2879), .B(net_2832), .A(net_2831) );
NOR2_X2 inst_3515 ( .A1(net_2397), .ZN(net_2346), .A2(net_1773) );
CLKBUF_X2 inst_10982 ( .A(net_10829), .Z(net_10830) );
CLKBUF_X2 inst_19112 ( .A(net_18959), .Z(net_18960) );
CLKBUF_X2 inst_13849 ( .A(net_11444), .Z(net_13697) );
INV_X2 inst_6332 ( .ZN(net_3025), .A(net_2988) );
SDFF_X2 inst_1270 ( .Q(net_7835), .D(net_7835), .SE(net_2730), .SI(net_2660), .CK(net_17030) );
CLKBUF_X2 inst_11593 ( .A(net_10127), .Z(net_11441) );
CLKBUF_X2 inst_12531 ( .A(net_12378), .Z(net_12379) );
AOI22_X2 inst_8001 ( .B1(net_8045), .A1(net_7841), .B2(net_6107), .ZN(net_6012), .A2(net_4400) );
NOR2_X2 inst_3448 ( .A2(net_3149), .ZN(net_2992), .A1(net_2991) );
INV_X4 inst_6088 ( .A(net_7249), .ZN(net_1959) );
CLKBUF_X2 inst_10123 ( .A(net_9543), .Z(net_9971) );
CLKBUF_X2 inst_16856 ( .A(net_16703), .Z(net_16704) );
CLKBUF_X2 inst_13032 ( .A(net_10114), .Z(net_12880) );
CLKBUF_X2 inst_14561 ( .A(net_14408), .Z(net_14409) );
INV_X4 inst_5361 ( .ZN(net_1143), .A(net_1142) );
CLKBUF_X2 inst_15602 ( .A(net_15449), .Z(net_15450) );
CLKBUF_X2 inst_12489 ( .A(net_12336), .Z(net_12337) );
CLKBUF_X2 inst_13049 ( .A(net_12896), .Z(net_12897) );
CLKBUF_X2 inst_15620 ( .A(net_15467), .Z(net_15468) );
SDFFR_X2 inst_2156 ( .Q(net_8274), .D(net_8274), .SI(net_3233), .SE(net_2996), .CK(net_18435), .RN(x6501) );
CLKBUF_X2 inst_18958 ( .A(net_12703), .Z(net_18806) );
CLKBUF_X2 inst_13389 ( .A(net_13145), .Z(net_13237) );
CLKBUF_X2 inst_12142 ( .A(net_11989), .Z(net_11990) );
CLKBUF_X2 inst_18411 ( .A(net_13987), .Z(net_18259) );
CLKBUF_X2 inst_19009 ( .A(net_18856), .Z(net_18857) );
INV_X4 inst_5417 ( .ZN(net_2570), .A(net_861) );
DFFR_X2 inst_7009 ( .QN(net_6314), .D(net_5793), .CK(net_14219), .RN(x6501) );
SDFFR_X2 inst_2515 ( .D(net_7367), .SE(net_2500), .SI(net_2499), .QN(net_231), .CK(net_16097), .RN(x6501) );
CLKBUF_X2 inst_17108 ( .A(net_16955), .Z(net_16956) );
CLKBUF_X2 inst_15798 ( .A(net_15645), .Z(net_15646) );
AOI222_X1 inst_8703 ( .A1(net_5031), .B2(net_5028), .C2(net_5027), .ZN(net_2788), .A2(net_2787), .B1(net_2786), .C1(net_1515) );
CLKBUF_X2 inst_12900 ( .A(net_11478), .Z(net_12748) );
XNOR2_X2 inst_117 ( .ZN(net_3173), .A(net_3039), .B(x2308) );
INV_X4 inst_5172 ( .ZN(net_3046), .A(net_2973) );
CLKBUF_X2 inst_13104 ( .A(net_12951), .Z(net_12952) );
CLKBUF_X2 inst_15195 ( .A(net_9363), .Z(net_15043) );
NAND2_X2 inst_4106 ( .ZN(net_5425), .A1(net_5239), .A2(net_5012) );
SDFF_X2 inst_465 ( .SI(net_8469), .Q(net_8469), .SE(net_3983), .D(net_3955), .CK(net_11022) );
SDFFR_X2 inst_2304 ( .D(net_3332), .SE(net_2313), .SI(net_431), .Q(net_431), .CK(net_16420), .RN(x6501) );
CLKBUF_X2 inst_11367 ( .A(net_9309), .Z(net_11215) );
CLKBUF_X2 inst_11701 ( .A(net_11548), .Z(net_11549) );
SDFFR_X2 inst_2173 ( .QN(net_7598), .SE(net_3144), .D(net_3128), .SI(net_1004), .CK(net_13503), .RN(x6501) );
DFFR_X2 inst_7048 ( .Q(net_7512), .D(net_4808), .CK(net_13741), .RN(x6501) );
OAI211_X2 inst_3214 ( .C1(net_1779), .ZN(net_1747), .B(net_1438), .A(net_783), .C2(net_205) );
CLKBUF_X2 inst_15039 ( .A(net_12103), .Z(net_14887) );
CLKBUF_X2 inst_16722 ( .A(net_13927), .Z(net_16570) );
SDFF_X2 inst_1905 ( .D(net_7268), .SI(net_7005), .Q(net_7005), .SE(net_6277), .CK(net_17050) );
CLKBUF_X2 inst_12940 ( .A(net_10346), .Z(net_12788) );
CLKBUF_X2 inst_11917 ( .A(net_11764), .Z(net_11765) );
CLKBUF_X2 inst_16201 ( .A(net_10570), .Z(net_16049) );
SDFFR_X2 inst_2264 ( .D(net_7390), .SE(net_2801), .SI(net_199), .Q(net_199), .CK(net_17770), .RN(x6501) );
CLKBUF_X2 inst_14925 ( .A(net_10523), .Z(net_14773) );
CLKBUF_X2 inst_18999 ( .A(net_18846), .Z(net_18847) );
CLKBUF_X2 inst_17163 ( .A(net_17010), .Z(net_17011) );
SDFFR_X1 inst_2697 ( .SI(net_7558), .SE(net_5043), .CK(net_12722), .RN(x6501), .Q(x3803), .D(x3803) );
XOR2_X2 inst_15 ( .Z(net_1451), .B(net_1450), .A(net_1333) );
CLKBUF_X2 inst_10196 ( .A(net_10043), .Z(net_10044) );
NAND4_X2 inst_3747 ( .ZN(net_4283), .A1(net_4033), .A2(net_4032), .A3(net_4031), .A4(net_4030) );
CLKBUF_X2 inst_11902 ( .A(net_9751), .Z(net_11750) );
NOR2_X2 inst_3496 ( .ZN(net_2162), .A1(net_1992), .A2(net_1874) );
CLKBUF_X2 inst_16025 ( .A(net_15872), .Z(net_15873) );
CLKBUF_X2 inst_13082 ( .A(net_12929), .Z(net_12930) );
CLKBUF_X2 inst_9830 ( .A(net_9166), .Z(net_9678) );
CLKBUF_X2 inst_13642 ( .A(net_13489), .Z(net_13490) );
SDFFR_X2 inst_2123 ( .SI(net_7186), .Q(net_7186), .D(net_6437), .SE(net_4362), .CK(net_17845), .RN(x6501) );
CLKBUF_X2 inst_12020 ( .A(net_11867), .Z(net_11868) );
MUX2_X2 inst_4918 ( .S(net_8901), .A(net_8252), .Z(net_5034), .B(net_1067) );
AOI222_X1 inst_8615 ( .ZN(net_5035), .A2(net_5034), .B1(net_5033), .A1(net_5031), .B2(net_5028), .C2(net_5027), .C1(net_1589) );
CLKBUF_X2 inst_17879 ( .A(net_17726), .Z(net_17727) );
CLKBUF_X2 inst_17736 ( .A(net_17583), .Z(net_17584) );
CLKBUF_X2 inst_14668 ( .A(net_13627), .Z(net_14516) );
CLKBUF_X2 inst_17110 ( .A(net_9703), .Z(net_16958) );
SDFF_X2 inst_349 ( .SI(net_8459), .Q(net_8459), .SE(net_3983), .D(net_3959), .CK(net_10047) );
CLKBUF_X2 inst_10690 ( .A(net_10537), .Z(net_10538) );
CLKBUF_X2 inst_14145 ( .A(net_11568), .Z(net_13993) );
CLKBUF_X2 inst_14381 ( .A(net_14228), .Z(net_14229) );
NAND2_X2 inst_4249 ( .A1(net_6907), .A2(net_5247), .ZN(net_5211) );
NAND2_X2 inst_4235 ( .A1(net_6900), .A2(net_5247), .ZN(net_5225) );
CLKBUF_X2 inst_13940 ( .A(net_9654), .Z(net_13788) );
CLKBUF_X2 inst_18967 ( .A(net_18814), .Z(net_18815) );
CLKBUF_X2 inst_17190 ( .A(net_12667), .Z(net_17038) );
CLKBUF_X2 inst_11507 ( .A(net_10226), .Z(net_11355) );
CLKBUF_X2 inst_13629 ( .A(net_12098), .Z(net_13477) );
CLKBUF_X2 inst_9570 ( .A(net_9417), .Z(net_9418) );
INV_X4 inst_6024 ( .A(net_7653), .ZN(net_508) );
CLKBUF_X2 inst_17030 ( .A(net_16877), .Z(net_16878) );
CLKBUF_X2 inst_14876 ( .A(net_14723), .Z(net_14724) );
CLKBUF_X2 inst_17965 ( .A(net_14338), .Z(net_17813) );
CLKBUF_X2 inst_17584 ( .A(net_17431), .Z(net_17432) );
CLKBUF_X2 inst_15725 ( .A(net_11247), .Z(net_15573) );
SDFFR_X2 inst_2252 ( .D(net_7393), .SE(net_2801), .SI(net_202), .Q(net_202), .CK(net_17775), .RN(x6501) );
CLKBUF_X2 inst_12289 ( .A(net_12136), .Z(net_12137) );
CLKBUF_X2 inst_12514 ( .A(net_12361), .Z(net_12362) );
CLKBUF_X2 inst_16095 ( .A(net_15942), .Z(net_15943) );
CLKBUF_X2 inst_17170 ( .A(net_9203), .Z(net_17018) );
NAND2_X2 inst_4229 ( .A1(net_6898), .A2(net_5247), .ZN(net_5231) );
CLKBUF_X2 inst_18253 ( .A(net_18100), .Z(net_18101) );
CLKBUF_X2 inst_12065 ( .A(net_11912), .Z(net_11913) );
SDFFR_X1 inst_2763 ( .QN(net_7568), .D(net_3981), .SE(net_3144), .SI(net_3110), .CK(net_13157), .RN(x6501) );
CLKBUF_X2 inst_10301 ( .A(net_10148), .Z(net_10149) );
CLKBUF_X2 inst_14334 ( .A(net_14181), .Z(net_14182) );
DFF_X1 inst_6798 ( .QN(net_8245), .D(net_4435), .CK(net_13586) );
CLKBUF_X2 inst_10554 ( .A(net_10401), .Z(net_10402) );
SDFF_X2 inst_761 ( .Q(net_8803), .D(net_8803), .SI(net_3954), .SE(net_3879), .CK(net_10526) );
NAND2_X2 inst_4867 ( .A1(net_8895), .ZN(net_1110), .A2(net_913) );
CLKBUF_X2 inst_13342 ( .A(net_10944), .Z(net_13190) );
OR3_X4 inst_2803 ( .A2(net_6113), .ZN(net_3003), .A1(net_1322), .A3(net_658) );
NAND2_X2 inst_4120 ( .ZN(net_5407), .A2(net_5230), .A1(net_5135) );
INV_X4 inst_5525 ( .ZN(net_666), .A(net_665) );
CLKBUF_X2 inst_9211 ( .A(net_9058), .Z(net_9059) );
INV_X4 inst_5097 ( .ZN(net_5696), .A(net_5669) );
CLKBUF_X2 inst_10003 ( .A(net_9566), .Z(net_9851) );
CLKBUF_X2 inst_16967 ( .A(net_16814), .Z(net_16815) );
SDFFR_X1 inst_2641 ( .D(net_6755), .SE(net_4506), .CK(net_9339), .RN(x6501), .SI(x2230), .Q(x2230) );
SDFF_X2 inst_1638 ( .Q(net_8154), .D(net_8154), .SI(net_2702), .SE(net_2538), .CK(net_18854) );
INV_X4 inst_5771 ( .A(net_9004), .ZN(net_845) );
CLKBUF_X2 inst_11450 ( .A(net_11297), .Z(net_11298) );
CLKBUF_X2 inst_17518 ( .A(net_17365), .Z(net_17366) );
CLKBUF_X2 inst_19062 ( .A(net_13999), .Z(net_18910) );
NOR4_X2 inst_3220 ( .ZN(net_2497), .A4(net_2496), .A2(net_2454), .A3(net_1072), .A1(net_848) );
CLKBUF_X2 inst_9812 ( .A(net_9104), .Z(net_9660) );
CLKBUF_X2 inst_18885 ( .A(net_18732), .Z(net_18733) );
AOI22_X2 inst_8177 ( .B1(net_8715), .A1(net_8493), .ZN(net_6077), .B2(net_4350), .A2(net_4349) );
INV_X4 inst_5354 ( .ZN(net_4320), .A(net_1802) );
CLKBUF_X2 inst_11983 ( .A(net_11830), .Z(net_11831) );
DFFR_X1 inst_7560 ( .Q(net_7642), .D(net_7633), .CK(net_15702), .RN(x6501) );
INV_X4 inst_5373 ( .ZN(net_1330), .A(net_1126) );
NAND2_X2 inst_4783 ( .ZN(net_1894), .A1(net_1570), .A2(net_1300) );
AND3_X2 inst_9047 ( .ZN(net_5275), .A2(net_4921), .A1(net_4701), .A3(net_4674) );
INV_X2 inst_6556 ( .A(net_7575), .ZN(net_3052) );
NAND4_X2 inst_3862 ( .ZN(net_1469), .A3(x2981), .A4(x2948), .A1(x2908), .A2(x2856) );
CLKBUF_X2 inst_17531 ( .A(net_17378), .Z(net_17379) );
INV_X2 inst_6532 ( .A(net_7492), .ZN(net_521) );
INV_X4 inst_5304 ( .ZN(net_2840), .A(net_2532) );
CLKBUF_X2 inst_10847 ( .A(net_10401), .Z(net_10695) );
CLKBUF_X2 inst_10482 ( .A(net_10329), .Z(net_10330) );
CLKBUF_X2 inst_14326 ( .A(net_14173), .Z(net_14174) );
SDFF_X2 inst_633 ( .SI(net_8547), .Q(net_8547), .SE(net_3979), .D(net_3953), .CK(net_10255) );
CLKBUF_X2 inst_18263 ( .A(net_18110), .Z(net_18111) );
CLKBUF_X2 inst_12837 ( .A(net_9619), .Z(net_12685) );
NAND2_X2 inst_4060 ( .ZN(net_5881), .A2(net_5766), .A1(net_3361) );
SDFFR_X2 inst_2285 ( .SI(net_7375), .SE(net_2793), .Q(net_234), .D(net_234), .CK(net_17828), .RN(x6501) );
CLKBUF_X2 inst_10500 ( .A(net_10347), .Z(net_10348) );
NAND2_X2 inst_4478 ( .A1(net_7163), .A2(net_4624), .ZN(net_4505) );
NOR2_X2 inst_3344 ( .ZN(net_5863), .A2(net_5713), .A1(net_2395) );
NOR2_X2 inst_3447 ( .ZN(net_3089), .A2(net_2961), .A1(net_1440) );
CLKBUF_X2 inst_11878 ( .A(net_11725), .Z(net_11726) );
CLKBUF_X2 inst_15968 ( .A(net_13118), .Z(net_15816) );
CLKBUF_X2 inst_17517 ( .A(net_17364), .Z(net_17365) );
DFFR_X2 inst_7199 ( .D(net_2373), .QN(net_223), .CK(net_14791), .RN(x6501) );
NAND2_X2 inst_4862 ( .A1(net_2807), .ZN(net_848), .A2(net_847) );
CLKBUF_X2 inst_19096 ( .A(net_18943), .Z(net_18944) );
NAND2_X2 inst_4663 ( .ZN(net_2218), .A1(net_2217), .A2(net_2216) );
CLKBUF_X2 inst_15220 ( .A(net_15067), .Z(net_15068) );
CLKBUF_X2 inst_10360 ( .A(net_10207), .Z(net_10208) );
SDFF_X2 inst_882 ( .Q(net_8561), .D(net_8561), .SI(net_3965), .SE(net_3878), .CK(net_12408) );
CLKBUF_X2 inst_13935 ( .A(net_9608), .Z(net_13783) );
CLKBUF_X2 inst_9848 ( .A(net_9695), .Z(net_9696) );
CLKBUF_X2 inst_13700 ( .A(net_13547), .Z(net_13548) );
OAI22_X2 inst_2938 ( .A1(net_2043), .ZN(net_2042), .B1(net_1857), .A2(net_1792), .B2(net_1136) );
AND2_X4 inst_9116 ( .A1(net_2827), .ZN(net_1506), .A2(net_1496) );
DFFS_X1 inst_6931 ( .D(net_6145), .CK(net_16354), .SN(x6501), .Q(x863) );
INV_X4 inst_5083 ( .ZN(net_5742), .A(net_5716) );
CLKBUF_X2 inst_15627 ( .A(net_15474), .Z(net_15475) );
CLKBUF_X2 inst_15802 ( .A(net_15649), .Z(net_15650) );
NAND2_X2 inst_4855 ( .A1(net_2810), .ZN(net_891), .A2(net_890) );
SDFF_X2 inst_1374 ( .Q(net_8188), .D(net_8188), .SI(net_2702), .SE(net_2561), .CK(net_18067) );
CLKBUF_X2 inst_17893 ( .A(net_9446), .Z(net_17741) );
SDFFR_X2 inst_2510 ( .Q(net_8996), .D(net_8996), .SI(net_2598), .SE(net_2562), .CK(net_17264), .RN(x6501) );
AND3_X4 inst_9046 ( .ZN(net_1819), .A1(net_1324), .A3(net_869), .A2(net_753) );
INV_X2 inst_6316 ( .ZN(net_3347), .A(net_3293) );
CLKBUF_X2 inst_15882 ( .A(net_11385), .Z(net_15730) );
CLKBUF_X2 inst_16532 ( .A(net_16379), .Z(net_16380) );
CLKBUF_X2 inst_19177 ( .A(net_9220), .Z(net_19025) );
CLKBUF_X2 inst_11548 ( .A(net_11395), .Z(net_11396) );
CLKBUF_X2 inst_14199 ( .A(net_14046), .Z(net_14047) );
CLKBUF_X2 inst_15184 ( .A(net_14052), .Z(net_15032) );
CLKBUF_X2 inst_16322 ( .A(net_16169), .Z(net_16170) );
DFF_X1 inst_6780 ( .Q(net_7558), .D(net_4592), .CK(net_10471) );
CLKBUF_X2 inst_18577 ( .A(net_10125), .Z(net_18425) );
NAND2_X2 inst_4398 ( .A1(net_7126), .A2(net_5166), .ZN(net_5059) );
NAND2_X2 inst_4165 ( .ZN(net_5347), .A2(net_5200), .A1(net_5090) );
SDFFR_X2 inst_2272 ( .SI(net_7383), .SE(net_2814), .Q(net_242), .D(net_242), .CK(net_17452), .RN(x6501) );
SDFF_X2 inst_1608 ( .Q(net_8145), .D(net_8145), .SI(net_2703), .SE(net_2541), .CK(net_14007) );
CLKBUF_X2 inst_11631 ( .A(net_11478), .Z(net_11479) );
SDFF_X2 inst_1484 ( .SI(net_7285), .Q(net_7062), .D(net_7062), .SE(net_6280), .CK(net_16213) );
SDFF_X2 inst_856 ( .SI(net_8638), .Q(net_8638), .D(net_3937), .SE(net_3885), .CK(net_11047) );
INV_X4 inst_5677 ( .A(net_7369), .ZN(net_1007) );
CLKBUF_X2 inst_18537 ( .A(net_16927), .Z(net_18385) );

endmodule
